��F6     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.5.1�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhN�verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ]�DhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��h3�f8�����R�(KhQNNNJ����J����K t�b�C              �?�t�bhUh'�scalar���hPC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hK�
node_count�M�nodes�h)h,K ��h.��R�(KM��h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h�hPK ��h�hPK��h�hPK��h�hbK��h�hbK ��h�hPK(��h�hbK0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@A         t                   �`@n�A��?L           ��@               Y       
             �?j?�]�?           `z@              :                    �?�	CO���?�            pt@                     	          ����?����l�?�            �p@        ������������������������       �        %             O@               #                   �n@(�Y7B��?�            `i@                                  �?��|Io��?P            �]@                                   �?և���X�?             @       	       
                   `j@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @               "                    �?�h����?L             \@                                 `_@���}<S�?2            @Q@        ������������������������       �                     2@                                  �_@�t����?%            �I@        ������������������������       �                      @                                  p`@Hm_!'1�?$            �H@                                   `@z�G�z�?             $@        ������������������������       �                     @                                   @K@����X�?             @       ������������������������       �                     @                                  @`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                      	          `ff�?�7��?            �C@        ������������������������       �                     �?                                  �_@P�Lt�<�?             C@       ������������������������       �                     ;@                                  pb@�C��2(�?             &@       ������������������������       �                     @                !                   `@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �E@        $       9                    �R@*�s���?4             U@       %       *       	          033�?^�pӵL�?3            @T@        &       '                   �p@z�G�z�?             $@        ������������������������       �                     @        (       )                   xs@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        +       .                    �?@�j;��?/            �Q@        ,       -       	             �?���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        /       2                    �?(;L]n�?(             N@        0       1                   `x@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        3       8                   �_@ �Jj�G�?$            �K@        4       5                    �?@4և���?	             ,@       ������������������������       �                     (@        6       7                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �D@        ������������������������       �                     @        ;       @                    �?�&�5y�?+             O@        <       =                   `X@z�G�z�?             $@        ������������������������       �                     �?        >       ?                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        A       T                   �c@D>�Q�?$             J@       B       C                     F@,���i�?            �D@        ������������������������       �                     �?        D       S                   p`@ףp=
�?             D@       E       N                    �L@�<ݚ�?             2@        F       M       	          ����?      �?             @       G       L       	          `ff�?���Q��?             @       H       I                    \@�q�q�?             @        ������������������������       �                     �?        J       K                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        O       P                    �?�8��8��?
             (@       ������������������������       �                     "@        Q       R                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        U       V                   @\@���|���?             &@        ������������������������       �                     @        W       X                    �P@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        Z       i                    �?�|R���??            �W@       [       b                   �c@     ��?,             P@        \       _                    [@"pc�
�?	             &@        ]       ^                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        `       a       	             п�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        c       d                   `a@���C��?#            �J@       ������������������������       �                     A@        e       f                    @L@�����?             3@       ������������������������       �                     $@        g       h                    ^@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        j       k                    ]@�P�*�?             ?@        ������������������������       �                     @        l       o                   �a@      �?             :@        m       n                   ps@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        p       q                    @M@������?             .@        ������������������������       �                      @        r       s                    �N@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        u       �                    �?�߸���?9            @        v       �       
             �?`�Q��?y            �e@       w       �                    �?�Ι����?A            @X@       x       y       
             �?h��Q(�?.            �P@        ������������������������       �                     &@        z       �                    �?      �?'             L@        {       ~                    �?     ��?             0@        |       }                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               �                    �?؇���X�?	             ,@        ������������������������       �                     @        �       �       	          @33�?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �       �                    @G@��Q���?             D@        �       �                   �n@      �?	             ,@       �       �                   �i@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          033�?8�Z$���?             :@       ������������������������       �        
             *@        �       �                   �c@�	j*D�?	             *@       �       �                    �?���|���?             &@        �       �                    b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �       	             @����X�?             @       �       �                    �N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     >@        �       �       	          ����?��
ц��?8            �S@       �       �                   �b@�	j*D�?$             J@        ������������������������       �                     1@        �       �                    �M@�xGZ���?            �A@       �       �                   �e@����"�?             =@        ������������������������       �                     @        �       �                    �? �o_��?             9@       �       �                   �b@�q�q�?             8@       �       �                   �i@�GN�z�?             6@        ������������������������       �                     �?        �       �                   �o@��s����?             5@        ������������������������       �                      @        �       �                    `@�	j*D�?             *@        �       �                   �c@z�G�z�?             @        ������������������������       �                     @        �       �                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   Pd@r�q��?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   c@�θ�?             :@       �       �                   �c@r�q��?             8@       ������������������������       �        
             .@        �       �       	          ����?X�<ݚ�?             "@       �       �                   �`@�q�q�?             @       �       �                    �?�q�q�?             @       �       �                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �K@ް� ��?�            t@       �       �                   �l@h��� �?�             n@        �       �                   �`@�|1)�?B            �Z@       �       �                   pa@`׀�:M�?2            �R@        �       �       
             �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        *            @P@        �       �                     B@      �?             @@        ������������������������       �                     �?        �       �                    @I@�g�y��?             ?@       ������������������������       �                     4@        �       �                    �?�C��2(�?             &@       ������������������������       �                      @        �       �       	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   Ph@L/)Lr��?L            �`@       �       �       
             �?\|/��j�?K            �`@        �       �                    �?H�z�G�?             D@        �       �                    �?      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        �       �                   �f@����X�?             <@       �       �                    �?z�G�z�?             9@       �       �                    �?r�q��?             8@        ������������������������       �                     @        ������������������������       �        
             4@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        5             W@        ������������������������       �                     @        �       �                   Pa@     ��?2             T@       �       �                    �?j���� �?             A@       �       �                   �a@J�8���?             =@        ������������������������       �                     @        �       �                   �a@R�}e�.�?             :@        ������������������������       �                     @        �       �                    �M@�q�q�?             5@       �       �       	          833�?z�G�z�?
             .@        �       �                    �?      �?              @       �       �                   (q@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   a@�q�q�?             @       �       �                   0b@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �m@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?�q��/��?             G@       �       �                    �?@4և���?             E@        ������������������������       �                     4@        �                         Ps@��2(&�?             6@       �       �                   �b@�����?             5@       ������������������������       �                     .@        �       �                   pk@�q�q�?             @        ������������������������       �                     �?        �              	          @33�?z�G�z�?             @       �       �                   `c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�b�values�h)h,K ��h.��R�(KMKK��hb�BP  >��=���?a�a��?��i�?�9K��?�a\&9�?��h���?үz�@�?���W��?              �?���/N�?Ztl��?:�:��?��O��O�?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?۶m۶m�?�$I�$I�?d!Y�B�?ӛ���7�?              �?�?<<<<<<�?      �?        9/���?Y�Cc�?�������?�������?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?�A�A�?��[��[�?      �?        (�����?���k(�?              �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?              �?z��y���?b�a��?�<ݚ�?���Hx�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        H���@��?w�'�K�?F]t�E�?]t�E]�?      �?                      �?�?�������?�������?�������?              �?      �?        ��)A��?k߰�k�?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?                      �?      �?        �1�c��?:�s�9�?�������?�������?              �?�q�q�?�q�q�?      �?                      �?vb'vb'�?b'vb'v�?8��18�?�����?      �?        �������?�������?�q�q�?9��8���?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?              �?      �?        &N��[��?�c�H;�?     ��?      �?F]t�E�?/�袋.�?      �?      �?      �?                      �?�q�q�?�q�q�?      �?                      �?\�琚`�?"5�x+��?      �?        Q^Cy��?^Cy�5�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�Zk����?�RJ)���?              �?      �?      �?/�袋.�?F]t�E�?      �?                      �?�?wwwwww�?              �?�$I�$I�?۶m۶m�?      �?                      �?�Zk����?SJ)��R�?{�G�z�?��(\���?���fy�?�Y�D�a�?z�rv��?�Wc"=P�?              �?      �?      �?      �?      �?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?F]t�E�?/�袋.�?              �?      �?        �������?333333�?      �?      �?ffffff�?333333�?              �?      �?                      �?;�;��?;�;��?              �?;�;��?vb'vb'�?F]t�E�?]t�E]�?      �?      �?      �?                      �?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?              �?              �?�;�;�?�؉�؉�?vb'vb'�?;�;��?      �?        �_�_�?�A�A�?	�=����?�i��F�?              �?
ףp=
�?�Q����?�������?�������?�袋.��?]t�E�?              �?z��y���?�a�a�?      �?        vb'vb'�?;�;��?�������?�������?              �?      �?      �?              �?      �?              �?                      �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        �؉�؉�?ى�؉��?UUUUUU�?�������?              �?�q�q�?r�q��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?      �?        J�#��?�rp�_��?�=&�=&�?�ξ?W�9�&�?"5�x+��?��L��?к����?�q�q�?�q�q�?              �?      �?              �?              �?      �?              �?��{���?�B!��?      �?        ]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?      �?                      �?e�+H��?n�Q�ߦ�?m��&�l�?N6�d�M�?333333�?ffffff�?      �?      �?      �?                      �?�$I�$I�?�m۶m��?�������?�������?UUUUUU�?�������?      �?                      �?      �?              �?              �?                      �?      �?      �?ZZZZZZ�?�������?|a���?�rO#,��?      �?        �;�;�?'vb'vb�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?333333�?�������?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?�������?�������?      �?                      �?�B����?��Mozӻ?n۶m۶�?�$I�$I�?      �?        ��.���?t�E]t�?=��<���?�a�a�?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ[�|/hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKͅ�h��B@3         �       
             �?��t�?O           ��@              Y                   �b@`U��Չ�?a           Ȁ@              .                    �?\Q�����?!           P{@                      	          @33�?��H�&p�?d            �b@                                   �F@XB���?&             M@                                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        	                           �? pƵHP�?!             J@       
                           �?XB���?             =@       ������������������������       �                     4@                                  �Z@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@                      	          ����?n�C���?>            �V@                                  �b@����"�?             =@                                 �m@�	j*D�?             :@                                  �?��.k���?             1@                                 @]@�	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @                                  `_@��a�n`�?)             O@        ������������������������       �                     5@               !       
             �?�p ��?            �D@                                  �`@���Q��?             @        ������������������������       �                     �?                                   `m@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        "       #                    �N@�����H�?             B@       ������������������������       �                     6@        $       )                   �`@����X�?
             ,@        %       &                    �?      �?             @        ������������������������       �                      @        '       (                   `^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        *       +                    �Q@ףp=
�?             $@       ������������������������       �                     @        ,       -                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        /       :                   �[@p�qG�?�             r@        0       9                    �O@���!pc�?            �@@       1       2                    �E@z�G�z�?             >@        ������������������������       �                      @        3       4       	          ����?���!pc�?             6@        ������������������������       �                     @        5       8                   �m@ҳ�wY;�?
             1@       6       7                   �]@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ;       F                   0`@�D�e���?�            �o@       <       A                    �?�o"Q9a�?r            �f@        =       @                   @_@$�q-�?             *@        >       ?                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        B       C                    �R@ �3_<�?k             e@       ������������������������       �        i            @d@        D       E                   �p@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        G       N                    �?@-�_ .�?5            �R@        H       M       	          033�?     ��?             0@       I       J       	             �?�z�G��?             $@        ������������������������       �                     @        K       L                   �a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        O       X       	          ����? _�@�Y�?)             M@        P       Q                    �?      �?             0@        ������������������������       �                     @        R       W                   0a@�����H�?             "@        S       T                   �a@�q�q�?             @        ������������������������       �                     �?        U       V                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     E@        Z       i                    �?4��@���?@             Y@        [       \                   Pc@�q�q�?            �C@        ������������������������       �                      @        ]       d                    �?�P�*�?             ?@        ^       c                   �e@������?             .@       _       b                   �c@�8��8��?             (@        `       a       	          `ff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        e       h       	             @      �?
             0@       f       g                    �?��S�ۿ?	             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     �?        j       k                   �Q@ҐϿ<��?(            �N@        ������������������������       �                     (@        l                          �f@և���X�?!            �H@       m       r                    �?F�����?            �F@        n       o                     K@      �?
             0@        ������������������������       �                      @        p       q                    @N@      �?              @        ������������������������       �                      @        ������������������������       �                     @        s       ~                    �?l��[B��?             =@       t       y                    �?���Q��?             9@        u       v                    @G@�����H�?             "@       ������������������������       �                     @        w       x                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        z       }                   �q@     ��?
             0@       {       |                   @d@      �?	             (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @E@
��`C2�?�            �w@        �       �                    �? \� ���?            �H@       �       �                    �Q@ܷ��?��?             =@       �       �       	          ����@4և���?             <@        ������������������������       �                     �?        �       �                   �`@ 7���B�?             ;@        �       �                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             2@        ������������������������       �                     �?        �       �                    �?�G�z��?             4@       �       �                    \@�	j*D�?             *@        ������������������������       �                     @        �       �                    �J@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �L@�#@���?�            �t@       �       �       	             @     >�?�             p@       �       �                    �?�j�}��?�            �o@        �       �                    �H@��P���?            �D@       �       �                   `\@և���X�?             5@        ������������������������       �                     @        �       �                    �?      �?             0@       ������������������������       �        	             (@        ������������������������       �                     @        ������������������������       �                     4@        �       �       	            �?��o�]�?�            �j@       �       �                    �?@t�!�a�?r            �f@       ������������������������       �        M             ^@        �       �                   c@0�z��?�?%             O@        �       �                   �b@ ��WV�?             :@       ������������������������       �                     9@        ������������������������       �                     �?        ������������������������       �                     B@        �       �                    �?      �?             @@        �       �                   0l@���Q��?             @        ������������������������       �                      @        �       �       	          pff�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @L@ 7���B�?             ;@       ������������������������       �                     :@        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          `ff�?�I�w�"�?1             S@       �       �                    �?���-T��?&             O@        �       �                    �?�E��ӭ�?             2@       �       �                   �b@     ��?             0@       ������������������������       �                     "@        �       �                   �_@և���X�?             @        ������������������������       �                     @        �       �                   �a@      �?             @        �       �                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    @M@�C��2(�?             F@        �       �                    �?      �?             @        �       �                   �q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   ht@P�Lt�<�?             C@       ������������������������       �                     B@        �       �                   �w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@X�Cc�?             ,@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        �       �                   @a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  |&�{&��?�l�l�?vH�w���?������?��c���?.�3j��?�IA��U�?��o�j�?�{a���?GX�i���?UUUUUU�?�������?      �?                      �?;�;��?'vb'vb�?�{a���?GX�i���?              �?�q�q�?�q�q�?      �?                      �?              �?���?�x��x��?	�=����?�i��F�?vb'vb'�?;�;��?�������?�?vb'vb'�?;�;��?              �?      �?                      �?      �?                      �?�c�1Ƹ?�s�9��?              �?��+Q��?Q��+Q�?�������?333333�?      �?              �?      �?              �?      �?        �q�q�?�q�q�?              �?�$I�$I�?�m۶m��?      �?      �?      �?              �?      �?              �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?t�E]t�?F]t�E�?�������?�������?              �?t�E]t�?F]t�E�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �???????�?�rS�<��?6��{��?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?              �?�a�ax?�<��<��?              �?UUUUUU�?�������?              �?      �?        к����?S�n0E�?      �?      �?333333�?ffffff�?              �?333333�?�������?      �?                      �?              �?�{a���?#,�4�r�?      �?      �?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?�G�z�?�(\����?UUUUUU�?UUUUUU�?      �?        �RJ)���?�Zk����?�?wwwwww�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?      �?�������?�?      �?                      �?              �?mާ�d�?������?              �?۶m۶m�?�$I�$I�?؂-؂-�?�>�>��?      �?      �?              �?      �?      �?      �?                      �?���=��?GX�i���?333333�?�������?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?                      �?      �?                      �?      �?        ��{��?�Ex^��?և���X�?
^N��)�?a���{�?��=���?�$I�$I�?n۶m۶�?      �?        h/�����?	�%����?�q�q�?�q�q�?      �?                      �?              �?      �?        �������?�������?vb'vb'�?;�;��?      �?        333333�?�������?              �?      �?                      �?�%���?GS��r�?      �?      �?>>>>>>�?�?������?�����?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?        YQ�@�?�Ե��?0��/���?h�h�v?      �?        |���{�?�B!��?O��N���?;�;��?      �?                      �?      �?              �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?	�%����?h/�����?      �?                      �?              �?����k�?�5��P�?[k���Z�?�RJ)���?�q�q�?r�q��?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?      �?                      �?              �?              �?]t�E�?F]t�E�?      �?      �?      �?      �?      �?                      �?      �?        ���k(�?(�����?      �?              �?      �?              �?      �?        �m۶m��?%I�$I��?              �?r�q��?�q�q�?              �?�������?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJh�rehG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�B         �                    �?Ly�'^��?L           ��@              _       
             �? �^���?f           ��@               B                   �`@m��1��?�             j@                                 0a@���)z�?N            �`@                                   Y@r�q��?             E@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        	       
                    �?�ݜ�?            �C@       ������������������������       �                     =@                      
             �?      �?             $@                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @                                  c@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                    D@���L��?5            �V@                                  @_@�<ݚ�?             "@                                  f@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?               %       	            �?�{��?.            �T@                                   �?R�}e�.�?             :@        ������������������������       �                     (@                                  �h@      �?             ,@        ������������������������       �                     @                       
             �?�z�G��?             $@        ������������������������       �                      @        !       $                    �F@      �?              @        "       #                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        &       3                    m@      �?             L@        '       2                    @M@���|���?             6@       (       1                    @      �?	             0@       )       *                    �F@�n_Y�K�?             *@        ������������������������       �                     �?        +       0                   l@�q�q�?             (@       ,       /                    �?�q�q�?             @       -       .       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        4       5                   �\@@�0�!��?             A@        ������������������������       �                     �?        6       A                     Q@6YE�t�?            �@@       7       @                    �?      �?             @@       8       ?                    �O@������?
             1@       9       >                    r@����X�?             ,@       :       =                    �?      �?              @       ;       <                    �K@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     �?        C       P                   �b@�7�QJW�?7            �R@       D       M       	          `ff@�>����?)             K@       E       J                    @`�q�0ܴ?$            �G@       F       I                   @]@ qP��B�?!            �E@       G       H                    �R@P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        ������������������������       �                     7@        K       L                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        N       O       
             �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        Q       \                    �N@և���X�?             5@       R       [                    �K@     ��?
             0@       S       X                    @      �?              @       T       W                   �c@z�G�z�?             @        U       V                    i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Y       Z                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ]       ^       	          ���@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        `       �       	          `ff @�ˠTX�?�             v@       a       r                   �]@� �ֺ��?�            pu@        b       m                    @L@��ga�=�?-            �P@       c       f                   �b@�:�B��?&            �M@       d       e                    ]@Pa�	�?            �@@       ������������������������       �                     @@        ������������������������       �                     �?        g       h                    �?$��m��?             :@        ������������������������       �                     @        i       j                   @m@�KM�]�?             3@       ������������������������       �                     &@        k       l                   @c@      �?              @        ������������������������       �                      @        ������������������������       �                     @        n       o       	             �?      �?              @        ������������������������       �                      @        p       q                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        s       z                   @E@Xe�&��?�            @q@        t       u                     K@      �?             0@        ������������������������       �                     @        v       w                   �a@���!pc�?	             &@       ������������������������       �                     @        x       y                    �P@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        {       |                   @i@����?�            @p@        ������������������������       �        .             S@        }       �                   �g@ �r�ѷ?t             g@       ~       �                    @L@ ��^og�?s            �f@              �       	          ����?�Ŗ�Pw�?Z            @a@       �       �                    �?`�߻�ɒ?I             [@        �       �                    �?P���Q�?             4@       �       �                    �?      �?             0@        ������������������������       �                     @        �       �                    �?$�q-�?             *@        ������������������������       �                     @        �       �                   �b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        =             V@        ������������������������       �                     >@        �       �       	          033�?���V��?            �F@       �       �                    @tk~X��?             B@       �       �                   pa@<���D�?            �@@        ������������������������       �        	             4@        �       �                     P@�	j*D�?	             *@       �       �                     N@      �?              @       �       �                    �L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?x疑��?�            `v@        �       �                    �?�7����?            �G@       �       �       
             �?�	j*D�?            �C@       �       �                    �J@����>�?            �B@        �       �                    �I@���Q��?             4@       �       �                    �?�t����?	             1@       �       �                    �C@�n_Y�K�?             *@        ������������������������       �                      @        �       �                   �k@�eP*L��?             &@        ������������������������       �                     @        �       �                   `c@����X�?             @       �       �                    @I@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@�t����?             1@        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �b@���%;��?�            ps@       �       �       
             �?4�Nx��?�            �q@       �       �                   �U@�Jƴ�o�?�            �o@        ������������������������       �                     �?        �       �                    �?h�����?�            �o@       �       �                    �L@�Ń��̧?�            @j@       �       �                   hp@Xc!J�ƴ?L            �]@       �       �                   �a@��S�ۿ?2            �R@       �       �                    �?x�}b~|�?'            �L@       �       �                   �_@�IєX�?"            �I@       �       �                    �?ףp=
�?             >@        ������������������������       �                     @        �       �                   �f@H%u��?             9@        ������������������������       �                     "@        �       �                     L@     ��?
             0@       �       �                    @K@@4և���?	             ,@       ������������������������       �                     &@        �       �       	          `ff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     5@        �       �                   �X@�q�q�?             @        ������������������������       �                     �?        �       �                   �^@z�G�z�?             @        ������������������������       �                      @        �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        ������������������������       �                    �E@        ������������������������       �        ;             W@        �       �                   �[@�����?             E@        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �N@�7��?            �C@       �       �                    n@�����?             5@       �       �                   �Q@�X�<ݺ?	             2@        �       �                     M@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �       	             �?�q�q�?             @        ������������������������       �                     �?        �       �                   0b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             2@        �       �                    �?�z�G��?             >@       �       �                   �q@r�q��?             8@       �       �       	             �?��2(&�?             6@        �       �                    n@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             0@        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �                          �?X�Cc�?             <@       �       �                    �K@z�G�z�?             4@       �       �       
             �?$�q-�?             *@        ������������������������       �                     @        �       �                    @I@�����H�?             "@        ������������������������       �                     @        �       �                   pf@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                 �d@և���X�?             @                                �?z�G�z�?             @                    	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                �l@      �?              @        ������������������������       �                     @        	      
      	          ���@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  ȫ�rV��?���T8�?B�A��?|�W|�W�?��؉���?;�;��?��9����?� れ�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?        �i�i�?\��[���?              �?      �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �����?�!�!�?�q�q�?9��8���?      �?      �?              �?      �?              �?        ��18�?������?�;�;�?'vb'vb�?              �?      �?      �?      �?        333333�?ffffff�?      �?              �?      �?      �?      �?              �?      �?                      �?      �?      �?]t�E]�?F]t�E�?      �?      �?ى�؉��?;�;��?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?              �?      �?              �?        ZZZZZZ�?�������?              �?'�l��&�?e�M6�d�?      �?      �?xxxxxx�?�?�m۶m��?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?              �?                      �?0��b�/�?t�@�t�?h/�����?�Kh/��?W�+�ɥ?��F}g��?�}A_З?��}A�?�������?ffffff�?              �?      �?                      �?      �?      �?              �?      �?        �$I�$I�?�m۶m��?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?      �?      �?�������?�������?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?                      �?F]t�E�?�E]tѽ?��U��?OZQ%�?��[���?�1���?�c+����?�pR���?|���?|���?      �?                      �?�N��N��?vb'vb'�?              �?�k(���?(�����?      �?              �?      �?              �?      �?              �?      �?      �?        UUUUUU�?�������?              �?      �?        `��k�?�%~F��?      �?      �?              �?F]t�E�?t�E]t�?      �?              �?      �?      �?                      �?Gn�Fn��?�����?      �?        �7��Mo�?��,d!�?��Z9��?�"Qj�a�?��?���?ہ�v`�}?B{	�%��?h/�����?ffffff�?�������?      �?      �?      �?        �؉�؉�?;�;��?      �?        �������?�������?      �?                      �?      �?              �?              �?        [�[��?�>�>��?r�q��?9��8���?|���?|���?      �?        vb'vb'�?;�;��?      �?      �?�������?�������?              �?      �?                      �?      �?                      �?      �?                      �?              �?59ȼ��?��fh�>�?G}g����?]AL� &�?;�;��?vb'vb'�?���L�?�u�)�Y�?�������?333333�?�������?�������?ى�؉��?;�;��?              �?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?              �?      �?        �?<<<<<<�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?              �?      �?        S���߷?V()��?��Ȇ�/�?��&���?�5g"�<�?��ٝ4��?      �?        �$I�$I�?�m۶m��?�a�a�?��<��<�?�pR�履?�؊���?�?�������?Lg1��t�?�YLg1�?�?�?�������?�������?              �?���Q��?)\���(�?              �?      �?      �?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?�a�a�?=��<���?UUUUUU�?UUUUUU�?              �?      �?        �A�A�?��[��[�?�a�a�?=��<���?�q�q�?��8��8�?      �?      �?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?333333�?ffffff�?UUUUUU�?�������?t�E]t�?��.���?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?�������?UUUUUU�?      �?                      �?�m۶m��?%I�$I��?�������?�������?;�;��?�؉�؉�?              �?�q�q�?�q�q�?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?�������?�������?      �?      �?              �?      �?                      �?      �?              �?      �?      �?        333333�?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ?PEhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�F         �       	          033�?�6𿸴�?G           ��@              C                    �K@����#�?9           �@                     
             �?������?�            @u@                      	          833�?��p �?0            �T@              
                    �?@4և���?"             L@               	                    �?�q�q�?             @                                  �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                                   g@`2U0*��?             I@                                 �`@@�E�x�?            �H@       ������������������������       �                     E@                                    F@؇���X�?             @                                  0a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                  �p@���B���?             :@                                 �Q@���}<S�?             7@                                   �I@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             1@        ������������������������       �                     @               B                   �f@�^龆��?�             p@              %                    P@     G�?�             p@               $                   `b@և���X�?             ,@              #                    �?z�G�z�?             $@              "                   �\@�����H�?             "@                !                     H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        &       3                    �?𯁷��?�            @n@        '       0       	          pff�?��2(&�?             F@       (       /                    @F@�˹�m��?             C@        )       *                   �d@     ��?             0@        ������������������������       �                      @        +       ,                    @E@@4և���?             ,@       ������������������������       �                     (@        -       .                    j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        1       2                     F@      �?             @        ������������������������       �                     @        ������������������������       �                     @        4       =                   �f@��		v�?}            �h@       5       6                   �b@@>ZAɥ�?u            `g@       ������������������������       �        >            @X@        7       8                   c@�X�<ݺ?7            �V@        ������������������������       �                      @        9       <                    �?�zvܰ?6             V@        :       ;                   �k@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        3            �T@        >       ?                    @C@"pc�
�?             &@       ������������������������       �                     @        @       A                   �f@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        D       _                   `_@�t��?k            �d@        E       X                    �?d}h���?-            �Q@       F       M       
             �?�7����?!            �G@       G       H       	          ����?XB���?             =@       ������������������������       �                     7@        I       L       	          hff�?r�q��?             @        J       K                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        N       O                   �`@�q�q�?             2@        ������������������������       �                      @        P       U                    �?���Q��?             $@        Q       R                    [@z�G�z�?             @        ������������������������       �                     @        S       T                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        V       W                   �]@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        Y       ^                   8r@���}<S�?             7@       Z       [                    �M@���7�?             6@       ������������������������       �                     2@        \       ]                   @V@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        `       q       
             �?�o+��?>            �W@        a       b                    `@�θ�?            �C@        ������������������������       �                     @        c       j                    �?r�q��?             B@       d       i                    �?���7�?             6@        e       h                    �?      �?             @       f       g                    c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     2@        k       p                   �c@X�Cc�?
             ,@       l       o                    �?"pc�
�?             &@       m       n                   �b@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        r       s                   �b@d}h���?$             L@        ������������������������       �                     8@        t                           �?      �?             @@        u       |       	          ����?�eP*L��?
             &@       v       w                    �L@      �?              @        ������������������������       �                     @        x       {                    �?z�G�z�?             @       y       z                   f@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        }       ~                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �c@����X�?             5@        �       �                    �?      �?              @       �       �                   @a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        �       �                   �c@:D?�H�?           �y@       �       �                    �R@R��+bH�?�            �v@       �       �                   �Q@�
d�<u�?�            0v@        ������������������������       �                      @        �       �                    �?�lY���?�            v@       �       �                    �J@ 
/'	�?�            pq@        �       �                   @X@��8����?<             X@        �       �       
             �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?ą%�E�?8            @V@       �       �                   �V@�G�V�e�?,             Q@        ������������������������       �                      @        �       �                   @e@��IF�E�?+            �P@        ������������������������       �                     &@        �       �                    �?X�;�^o�?&            �K@        ������������������������       �                      @        �       �                    �?��0{9�?             �G@       �       �                   `b@ףp=
�?             D@       �       �                    �H@�IєX�?             A@       ������������������������       �                     6@        �       �       	             �?r�q��?	             (@       �       �                    �I@����X�?             @       �       �                   �]@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    ]@և���X�?             @        ������������������������       �                      @        �       �                     H@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        �       �                    c@ �ղ?y            �f@       �       �                    �?�O���h�?w            �f@        �       �                    ]@؇���X�?             5@        �       �                   �R@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �`@�IєX�?
             1@        �       �       	             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                   �_@Уp=
ע?j             d@        �       �                    I@ �#�Ѵ�?             �E@        �       �                   `_@؇���X�?             ,@       �       �                    �?$�q-�?
             *@        �       �                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     =@        �       �       	          ����?�6H�Z�?J            @]@        �       �                    �K@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �        >            �W@        �       �                   c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �e@�r*e���?2            �R@       �       �                   �`@L�w�=�?0            �Q@       �       �                     P@z�G�z�?             D@       �       �                   �c@     ��?             @@       �       �                    �?��S�ۿ?             >@        �       �       	          033�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @M@ 7���B�?             ;@       ������������������������       �        
             1@        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                   P`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                      @        �       �                    @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          `ff�?��S���?             >@        �       �                   �f@�θ�?             *@        ������������������������       �                      @        �       �                   @b@�C��2(�?             &@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@ҳ�wY;�?             1@        ������������������������       �                      @        �       �       
             �?������?             .@       �       �       	          `ff�?r�q��?             (@        �       �       	          `ff�?�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �                         �d@����3��?#             J@        �                          �?�q�q�?             8@       �                         �q@�����?             5@                                 �?�X�<ݺ?             2@       ������������������������       �                     ,@                                 �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?                    	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        	                         �?      �?             <@       
                        �e@���|���?             6@                    	          ���@���Q��?             $@                               e@և���X�?             @        ������������������������       �                     @                                Pe@      �?             @        ������������������������       �                      @                                 b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  I@r�q��?             (@                                �?�C��2(�?             &@       ������������������������       �                     "@                                �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KMKK��hb�B�  (Dҵ��?l�����?;�����?�'�ɂn�?xxxxxx�?�?��18��?>�cp>�?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?{�G�z�?���Q��?9/���?և���X�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��؉���?ى�؉��?ӛ���7�?d!Y�B�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?I[Җ�%�?�%mI[Ҷ?     `�?      �?۶m۶m�?�$I�$I�?�������?�������?�q�q�?�q�q�?      �?      �?      �?                      �?              �?      �?              �?        �
�G�?j�V���?��.���?t�E]t�?��P^Cy�?^Cy�5�?      �?      �?              �?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?              �?              �?      �?      �?                      �?�y;Cb��?ogH���?%��j�$�?a�2a�?      �?        ��8��8�?�q�q�?              �?颋.���?t�E]t�?�������?333333�?      �?                      �?      �?        /�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?`�1`�?�r�,���?۶m۶m�?I�$I�$�?G}g����?]AL� &�?�{a���?GX�i���?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?333333�?�������?�������?              �?      �?      �?      �?                      �?333333�?�������?      �?                      �?d!Y�B�?ӛ���7�?F]t�E�?�.�袋�?              �?      �?      �?              �?      �?              �?        �+F��?�ĩ�sK�?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?F]t�E�?�.�袋�?      �?      �?      �?      �?      �?                      �?              �?              �?�m۶m��?%I�$I��?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        I�$I�$�?۶m۶m�?      �?              �?      �?]t�E�?t�E]t�?      �?      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �³��?�SB�?#����%�?w����6�?���3��?B�E��?      �?        �v���
�?D���G��?�gI��Y�?
���´�?UUUUUU�?�������?�$I�$I�?۶m۶m�?              �?      �?        ��g<�?�as���?�������?�������?      �?        '�l��&�?�l��&��?              �?J��yJ�?�־a��?              �?L� &W�?m�w6�;�?�������?�������?�?�?              �?UUUUUU�?�������?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?              �?��ݮ��?�/���?������?�0&q��?�$I�$I�?۶m۶m�?      �?      �?              �?      �?        �?�?�������?�������?      �?                      �?              �?333333�?ffffff�?�}A_Ч?�/����?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?���?�������?d!Y�B�?�Mozӛ�?      �?                      �?              �?      �?      �?              �?      �?        �u�)�Y�?0E>�S�?uPuP�?�W|�W|�?ffffff�?ffffff�?      �?      �?�?�������?UUUUUU�?UUUUUU�?              �?      �?        h/�����?	�%����?              �?�������?�������?              �?�������?�������?      �?                      �?      �?      �?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?�������?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?      �?              �?      �?      �?              �?      �?              �?      �?        �������?�������?      �?        �?wwwwww�?UUUUUU�?�������?UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        �������?UUUUUU�?      �?                      �?��N��N�?'vb'vb�?UUUUUU�?�������?=��<���?�a�a�?��8��8�?�q�q�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?]t�E]�?F]t�E�?�������?333333�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?              �?      �?                      �?�������?UUUUUU�?]t�E�?F]t�E�?      �?              �?      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�#jThG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�A         �       
             �?Np�����?C           ��@              #                    �?$���-�??           P~@               "                    �?      �?5            �S@                                  �?     x�?-             P@                                  �D@��P���?            �D@        ������������������������       �                      @                                  �\@:�&���?            �C@        ������������������������       �                     @        	                          hq@�#-���?            �A@       
                          �b@`Jj��?             ?@       ������������������������       �                     =@        ������������������������       �                      @                                  �q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                      	          ����?8����?             7@        ������������������������       �                     @                                   �?p�ݯ��?             3@                                 �o@     ��?             0@                      	             �?�q�q�?             @        ������������������������       �                      @                                    I@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   �?ףp=
�?             $@        ������������������������       �                     @                                   `@r�q��?             @                                  pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                !                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        $       k                    a@H߾���?
           py@       %       P                   �\@l������?�            �r@        &       E                    �?0�й���?X            @b@       '       >       	             @�IєX�?I            �]@       (       7                   `[@h㱪��?C            �[@       )       2                    �O@`���i��?6             V@       *       1                   @X@ ��PUp�?+            �Q@        +       ,                    �?(;L]n�?             >@        ������������������������       �                     ,@        -       .                   �W@      �?             0@       ������������������������       �        	             (@        /       0                     L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �D@        3       6                     P@�IєX�?             1@        4       5                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        8       9                   0l@�C��2(�?             6@        ������������������������       �                     (@        :       =                   �c@z�G�z�?             $@       ;       <                   �n@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ?       @                   Pn@�q�q�?             "@        ������������������������       �                     @        A       B                   �Z@      �?             @        ������������������������       �                     �?        C       D                     M@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        F       G                    �?�5��?             ;@        ������������������������       �                     "@        H       I       
             �?�����H�?             2@        ������������������������       �                     @        J       O                    �?r�q��?
             (@        K       N                   `Z@�q�q�?             @       L       M                   �^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Q       h                    @p�|�i�?e             c@       R       a                   P`@(;L]n�?c            �b@        S       `       	          ����?l�b�G��?+            �L@       T       _                   �r@<���D�?            �@@       U       \                    �?`Jj��?             ?@       V       W                    �?h�����?             <@        ������������������������       �                     @        X       Y       	          `ff�?���N8�?             5@       ������������������������       �                     3@        Z       [       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        b       g                     E@�L��ȕ?8            @W@        c       d                    b@      �?             @        ������������������������       �                      @        e       f                   `U@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        5            @V@        i       j                   @]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        l       �                    �J@ ��?�?M            @[@        m       �                   `o@nM`����?!             G@       n                          �m@��.k���?             A@       o       z                   �^@����"�?             =@        p       q                   pa@      �?
             0@        ������������������������       �                     @        r       u       	             �?�θ�?	             *@        s       t                    �H@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        v       w       	          033@ףp=
�?             $@       ������������������������       �                      @        x       y                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        {       ~                   ``@$�q-�?             *@        |       }                    @J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?�8��8��?	             (@       ������������������������       �                     @        �       �                   `]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?؇���X�?,            �O@        �       �                   �e@���7�?             6@       ������������������������       �                     4@        �       �                     N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?� ��1�?            �D@       �       �                   �`@     ��?             @@       ������������������������       �                     2@        �       �                   `l@d}h���?             ,@       �       �                    �?�����H�?             "@       �       �                    i@؇���X�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	             @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          `ff�?X�<ݚ�?             "@        ������������������������       �                      @        �       �                   �_@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@P@㞲��?           {@       �       �       	          ����?�3��j�?�            Ps@       �       �       	          ���ٿP#aE�?�            �p@        �       �                    @F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          833�? �q�q�?�            �p@       �       �                    �?г�wY;�?�            �m@        �       �                   @E@fP*L��?             F@        ������������������������       �                      @        �       �                    �?���H��?             E@        ������������������������       �                     "@        �       �                    ]@6YE�t�?            �@@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�8��8��?             8@       �       �                   �e@���N8�?             5@       ������������������������       �                     3@        �       �                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        n            @h@        �       �                    �E@8�Z$���?             :@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���7�?             6@        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        �       �                   `T@�lg����?            �E@        ������������������������       �                     (@        �       �                   �d@��� ��?             ?@       �       �                    �?�nkK�?             7@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     3@        �       �                   �e@      �?              @        �       �                    �G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?f���M�?F             _@        �       �                   �b@�����H�?             ;@        ������������������������       �                      @        �       �                    �?�S����?
             3@       �       �                   ps@�z�G��?             $@        ������������������������       �                     @        �       �                   @a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?lG:<�?7            @X@       �       �                   �r@�E��
��?             J@       �       �                   �]@(옄��?             G@        ������������������������       �                     $@        �       �                    �?�q�q�?             B@       �       �                    �?      �?             <@        �       �                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �X@r�q��?             8@        �       �                   �_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    b@P���Q�?
             4@       ������������������������       �                     ,@        �       �                   �b@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�<ݚ�?            �F@        �       �                    �?���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    ]@z�G�z�?             D@        ������������������������       �                     �?        �                         Ps@:�&���?            �C@       �       �                   Hp@$G$n��?            �B@       �       �                    @ףp=
�?             >@       �       �                    �Q@���7�?             6@       ������������������������       �        
             2@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @N@      �?              @        ������������������������       �                      @        ������������������������       �                     @                                 �a@����X�?             @                               @a@r�q��?             @        ������������������������       �                     @                                @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�Bp  ______�?PPPPPP�?�M��}�?��E̹ �?      �?      �?     ��?      �?������?�����?              �?�A�A�?�o��o��?              �?�A�A�?_�_�?���{��?�B!��?      �?                      �?      �?      �?              �?      �?        8��Moz�?d!Y�B�?              �?Cy�5��?^Cy�5�?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�k�s�?������?��c.��?+�3�=l�?����Ǐ�?����?�?�?��)A��?־a���?F]t�E�?F]t�E�?��V،?��ۥ���?�?�������?              �?      �?      �?              �?      �?      �?              �?      �?                      �?�?�?      �?      �?              �?      �?                      �?F]t�E�?]t�E�?              �?�������?�������?�q�q�?�q�q�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?333333�?�������?      �?                      �?/�����?h/�����?      �?        �q�q�?�q�q�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?^Cy�5�?�k(����?�?�������?p�}��?�Gp��?|���?|���?�B!��?���{��?�$I�$I�?�m۶m��?              �?�a�a�?��y��y�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?X`��?��~���?      �?      �?              �?      �?      �?              �?      �?                      �?      �?      �?              �?      �?        ���]8��?߅���]�?zӛ����?C���,�?�?�������?�i��F�?	�=����?      �?      �?              �?ى�؉��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?              �?      �?      �?                      �?;�;��?�؉�؉�?UUUUUU�?�������?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?�$I�$I�?۶m۶m�?F]t�E�?�.�袋�?              �?      �?      �?      �?                      �?������?������?      �?      �?              �?۶m۶m�?I�$I�$�?�q�q�?�q�q�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?              �?�������?333333�?      �?                      �?r�q��?�q�q�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        #Up�ѭ�?t�>v�H�?Z�Ϯ�?.�
��2�?�蛣o��?�qA��?      �?      �?      �?                      �?�������?UUUUUU�?�?�?颋.���?]t�E]�?              �?�0�0�?��y��y�?      �?        '�l��&�?e�M6�d�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?��y��y�?�a�a�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ;�;��?;�;��?      �?      �?              �?      �?        �.�袋�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?        }A_��?�}A_��?              �?�{����?�B!��?�Mozӛ�?d!Y�B�?      �?      �?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?      �?        ��RJ)��?��Zk���?�q�q�?�q�q�?      �?        (������?^Cy�5�?ffffff�?333333�?      �?              �?      �?              �?      �?              �?        ���fy�?���$2�?��؉���?;�;��?ӛ���7�?���,d�?              �?�������?�������?      �?      �?      �?      �?              �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?ffffff�?�������?      �?        �������?UUUUUU�?              �?      �?                      �?              �?9��8���?�q�q�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?              �?�A�A�?�o��o��?к����?���L�?�������?�������?�.�袋�?F]t�E�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?        �m۶m��?�$I�$I�?�������?UUUUUU�?      �?              �?      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�JvhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@D         �       	          ����?�6𿸴�??           ��@               /                   `@X�C��?            |@                                   �?�n_Y�K�?M            @]@                                   �?�r����?
             .@                      
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        	       *                    �?�\�u��?C            �Y@       
                          b@�Jhu4��?1            @R@                                   �?��a�n`�?             ?@                     	          @33�?`2U0*��?             9@                                 @b@�}�+r��?             3@       ������������������������       �                     1@                                  e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   \@�q�q�?             @        ������������������������       �                      @                      
             �?      �?             @                                 @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                  �[@X�Cc�?             E@                                   �?�X�<ݺ?             2@       ������������������������       �                      @                                   �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@                %                   `q@�q�q�?             8@       !       $       
             �?�����?             3@       "       #                   �_@�r����?	             .@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        &       )                    �J@z�G�z�?             @       '       (       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        +       ,                    �? 	��p�?             =@       ������������������������       �                     4@        -       .                     G@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        0       e                    �?�E���?�            �t@        1       V                    �L@�Q����?B            @\@       2       Q                    �?<�\`*��?1             U@       3       B                   �_@:-�.A�?&            �P@        4       ;                    ]@      �?             8@        5       6                   `i@�q�q�?             "@        ������������������������       �                      @        7       8                    �?؇���X�?             @        ������������������������       �                      @        9       :                    �H@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        <       =                    �?z�G�z�?             .@        ������������������������       �                     �?        >       ?                    �K@؇���X�?             ,@       ������������������������       �                     $@        @       A                    b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        C       D                    P@�ʈD��?            �E@        ������������������������       �                     �?        E       P                   �b@@4և���?             E@       F       G                   �b@������?            �D@        ������������������������       �        	             2@        H       K                    `@���}<S�?             7@        I       J                    d@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        L       O                   c@�IєX�?
             1@        M       N       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     �?        R       S                   ``@j���� �?             1@       ������������������������       �                      @        T       U                   �a@�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                      @        W       Z                    �?V�a�� �?             =@        X       Y                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        [       d                    �?8�Z$���?             :@       \       _                    �M@�	j*D�?             *@        ]       ^                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        `       c                   �^@z�G�z�?             $@        a       b                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        f       �                   �z@���qh�?�            @k@       g       z       
             �?<�*/�{�?�             k@        h       u                   Po@h+�v:�?             A@       i       l                   �_@����X�?             <@        j       k                   @W@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        m       p                    @G@p�ݯ��?
             3@        n       o                    @B@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        q       t                   �`@���Q��?             $@       r       s                    f@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        v       y                    �?r�q��?             @        w       x                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        {       |                    @L@��v$���?r            �f@       ������������������������       �        ]            �b@        }       ~                    �?     ��?             @@        ������������������������       �                     &@               �                    �?؇���X�?             5@       �       �                    �?�z�G��?             $@        �       �                    �?�q�q�?             @       �       �                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �?���Lr��?(           `}@        �       �       
             �?��6���?5             U@       �       �                    �?�u���?'            �N@       �       �                    _@:�&���?            �C@        �       �                   �n@      �?              @        �       �                   �Z@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @L@��a�n`�?             ?@        ������������������������       �                     (@        �       �                   hu@�S����?
             3@       �       �       
             �?�IєX�?	             1@        ������������������������       �                     @        �       �                    �?$�q-�?             *@        �       �                   �p@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        �       �       	          ����?�GN�z�?             6@        �       �                    @      �?              @       �       �       	          ����?����X�?             @       �       �                    @M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   @Z@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        �       �                   �b@���[�A�?�             x@       �       �       	          ���@`Er�ٍ�?�            �t@       �       �                   �`@��Fi�1�?�            0p@       �       �       	             �?����H�?z            `h@        �       �       
             �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                   �z@�f����?v             g@       �       �       	          pff�?��GEI_�?t            �f@       �       �                   �j@     p�?Q             `@       �       �                    �L@      �?-             R@        �       �                    @L@�'�`d�?            �@@       �       �                    �?$�q-�?             :@       �       �                    d@      �?             0@        ������������������������       �                      @        �       �       
             �?      �?              @       �       �                     E@؇���X�?             @        �       �                    b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   `@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?�7��?            �C@       �       �                   �X@������?             B@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     >@        �       �                   �c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �s@�h����?$             L@       ������������������������       �        !            �I@        �       �                    [@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �R@h㱪��?#            �K@       ������������������������       �        "            �J@        ������������������������       �                      @        �       �                   @X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �[@     ��?&             P@        ������������������������       �                      @        �       �       
             �?�>4և��?#             L@       �       �                    �? ���J��?            �C@        �       �       	          033@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     =@        �       �                   pb@��.k���?
             1@       �       �                    �?և���X�?             ,@       �       �                    @N@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @P�Lt�<�?-             S@       ������������������������       �        +             R@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �       	          ����?Np�����?&            �I@        �       �                   �d@�r����?             .@        ������������������������       �                     @        �       �                    �G@z�G�z�?             $@       ������������������������       �                     @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       
                  (p@*O���?             B@                                �]@D�n�3�?             3@        ������������������������       �                      @                                 �?ҳ�wY;�?             1@                    	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @              	                   `@r�q��?
             (@                    	          ���@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                @_@�t����?
             1@        ������������������������       �                      @                                0s@�<ݚ�?             "@                               �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�B  (Dҵ��?l�����?۶m۶��?I�$I�$�?ى�؉��?;�;��?�������?�?      �?      �?              �?      �?              �?        �?�������?ҤI�&M�?�-[�l��?�c�1Ƹ?�s�9��?{�G�z�?���Q��?(�����?�5��P�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        %I�$I��?�m۶m��?��8��8�?�q�q�?      �?        �������?�������?              �?      �?        �������?�������?^Cy�5�?Q^Cy��?�?�������?              �?      �?              �?        �������?�������?      �?      �?              �?      �?              �?        �{a���?������?              �?�q�q�?9��8���?      �?                      �?5QeWMT�?+�j�ʮ�?�c�:F�?�8�1�s�?=��<���?�a�a�?���@���?��~5&�?      �?      �?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?�������?�������?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?A_���?�}A_з?              �?n۶m۶�?�$I�$I�?p>�cp�?������?      �?        ӛ���7�?d!Y�B�?�������?UUUUUU�?      �?                      �?�?�?      �?      �?              �?      �?              �?                      �?ZZZZZZ�?�������?              �?9��8���?�q�q�?      �?                      �?a���{�?��{a�?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?;�;��?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?ش�,��?j?Y���?��G���?��K�%�?�������?xxxxxx�?�m۶m��?�$I�$I�?�q�q�?�q�q�?              �?      �?        ^Cy�5�?Cy�5��?�q�q�?�q�q�?              �?      �?        �������?333333�?�$I�$I�?۶m۶m�?              �?      �?              �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?.�u�y�?;ڼOqɐ?      �?              �?      �?      �?        ۶m۶m�?�$I�$I�?ffffff�?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �m۶m��?�$I�$I�?              �?      �?              �?                      �?�"��i�?I�>���?b�a��?=��<���?XG��).�?T\2�h�?�o��o��?�A�A�?      �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?�c�1Ƹ?�s�9��?              �?^Cy�5�?(������?�?�?              �?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?        �袋.��?]t�E�?      �?      �?�$I�$I�?�m۶m��?�������?�������?              �?      �?              �?      �?              �?      �?              �?              �?        �Mozӛ�?d!Y�B�?              �?      �?        ko��@��?%�T�/��?�X����?^�ti���?�Q:���?ʼk1���?PP�?��_��_�?333333�?ffffff�?      �?                      �?���;��?��X��?;ڼOqɰ?�d����?      �?     ��?      �?      �?'�l��&�?6�d�M6�?;�;��?�؉�؉�?      �?      �?              �?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�m۶m��?�$I�$I�?      �?                      �?�A�A�?��[��[�?�q�q�?�q�q�?UUUUUU�?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?        ��)A��?־a���?              �?      �?              �?      �?      �?                      �?      �?      �?      �?        �m۶m��?�$I�$I�?�A�A�?��-��-�?�������?�������?              �?      �?                      �?�������?�?۶m۶m�?�$I�$I�?      �?      �?      �?      �?              �?      �?                      �?�������?UUUUUU�?      �?                      �?      �?        (�����?���k(�?              �?      �?      �?      �?                      �?PPPPPP�?______�?�������?�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�q�q�?�q�q�?l(�����?(������?              �?�������?�������?�������?�������?      �?                      �?�������?UUUUUU�?333333�?�������?      �?                      �?      �?        �?<<<<<<�?              �?�q�q�?9��8���?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���GhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�G         �                    �?n�A��?C           ��@              !                   @E@hW����?4           @~@                      	          033�?�-���e�?P            �_@              	                    Z@ rpa�?;            @W@                      	          ���ܿ����X�?             @        ������������������������       �                      @                                  �X@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        
                          �b@��+��<�?7            �U@                                  �?�e���@�?2            @S@       ������������������������       �        "            �J@                      
             �? �q�q�?             8@       ������������������������       �                     1@                                   @M@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                      	          ����?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @                                  �U@"pc�
�?            �@@        ������������������������       �                      @                                   �?��� ��?             ?@       ������������������������       �                     4@                                  p`@���|���?             &@                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                      
             �?؇���X�?             @       ������������������������       �                     @                                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        "                          �a@��=����?�            `v@       #       R                    �?�[�|Tc�?�            �o@        $       9                   �l@�	#i���?E            �Z@        %       4       	          033�?�<ݚ�?!            �F@       &       '                    �?8�Z$���?            �C@        ������������������������       �                      @        (       -                   �b@�n`���?             ?@       )       ,       
             �?ȵHPS!�?             :@        *       +                   �_@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        .       3                   @`@���Q��?             @       /       0       
             �?      �?             @        ������������������������       �                      @        1       2                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        5       6       	          ����?�q�q�?             @        ������������������������       �                     @        7       8                   @^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        :       G       
             �?`՟�G��?$             O@       ;       B                    �?�q�q�?            �@@        <       A       	          `ff@�q�q�?             (@       =       >       	          ����?z�G�z�?             $@        ������������������������       �                     �?        ?       @                   �\@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        C       D                     M@؇���X�?             5@       ������������������������       �                     .@        E       F                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     @        H       I                   �b@�f7�z�?             =@        ������������������������       �                     @        J       K                    �I@�eP*L��?             6@        ������������������������       �                     @        L       M                   �_@�t����?             1@        ������������������������       �                     $@        N       Q                    �?����X�?             @       O       P                   �s@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        S       x       
             �?^	����?X            @b@       T       q                   @b@X��Oԣ�?M             _@       U       j                    �O@ >�֕�?B            @Z@       V       i                    �L@��8�$>�?;            @X@       W       h                   pp@F��}��?+            @R@       X       g                   �o@dP-���?            �G@       Y       `                   `_@���.�6�?             G@       Z       [                   @l@XB���?             =@       ������������������������       �                     3@        \       _                    \@ףp=
�?             $@        ]       ^       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        a       f       	          ����?�t����?
             1@       b       e                    �?r�q��?             (@        c       d                    ^@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@        ������������������������       �                     8@        k       l                   �Y@      �?              @        ������������������������       �                     @        m       n                    _@���Q��?             @        ������������������������       �                      @        o       p                    [@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        r       u                    a@D�n�3�?             3@       s       t       	          ���@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        v       w                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        y       z                    _@�X����?             6@        ������������������������       �                     @        {       |                   �`@b�2�tk�?	             2@        ������������������������       �                     @        }       ~                   pf@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   `f@T>D5j�?G            @Z@       �       �                    y@�8��8N�?A             X@       �       �                   �b@8v�YeK�?@            �W@        ������������������������       �                     ?@        �       �       
             �?     ��?+             P@       �       �                    �R@�O4R���?#            �J@       ������������������������       �        "             J@        ������������������������       �                     �?        �       �       	          033�?�eP*L��?             &@       �       �                   po@�q�q�?             "@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                     L@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        �       �       
             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?�HcJ]�?            {@        �       �                   �b@�fp�I��?i             d@       �       �       	          @33�?4A�,��?F            �Y@        �       �                    �?`2U0*��?             9@        �       �                   �_@r�q��?             @       ������������������������       �                     @        �       �                     C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        �       �                   �`@^Gث3��?4            �S@       �       �                    @P@؇���X�?            �A@       �       �                    @M@ 7���B�?             ;@        ������������������������       �                     (@        �       �                    �?��S�ۿ?             .@       �       �       	          ����?ףp=
�?             $@        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?              @        �       �                   @]@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?�K��&�?            �E@        ������������������������       �                     @        �       �       	             @�99lMt�?            �C@       �       �                   o@4���C�?            �@@       �       �                    �L@�q�q�?             2@       �       �                    �?      �?             $@       �       �                     H@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �[@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `P@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �b@�r����?             .@       ������������������������       �                     $@        �       �                    ]@���Q��?             @        ������������������������       �                     �?        �       �                   @q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �d@����S��?#             M@        �       �       	          `ff@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ���@�c�����?            �J@       �       �                    �?z�G�z�?             I@        �       �       	          `ff�?���N8�?             5@       �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                   d@      �?             @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �       �       
             �?8^s]e�?             =@        ������������������������       �                     @        �       �                   ``@$��m��?             :@       �       �                   pe@      �?	             0@       ������������������������       �                     $@        �       �                    @I@r�q��?             @       �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @z�G�z�?             $@        ������������������������       �                     @        �       �                   �c@      �?             @        ������������������������       �                     �?        �       �                   @b@�q�q�?             @        ������������������������       �                     �?        �       �                   e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                           R@0�>���?�            q@       �                          �?�f��'�?�            �p@        �       �                    c@0��_��?            �J@       �       �                    �L@ "��u�?             I@       �       �                    @G@�?�|�?            �B@        ������������������������       �                     5@        �       �                    �?      �?	             0@       ������������������������       �                     $@        �       �                   �]@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ��� @8�Z$���?
             *@       �       �                    �?�8��8��?	             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �       �                   `c@�q�q�?             @        ������������������������       �                     �?        �                            @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 ]@���*}ǫ?�            �j@                                 �?ףp=
�?             >@       ������������������������       �                     1@                                �V@�θ�?             *@        ������������������������       �                     �?                                `m@r�q��?             (@       ������������������������       �                     @        	      
                  �n@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                 �?�x�V�?r             g@                               �c@����7�?k             f@                   	            �?`�E���?=            @X@                                t@ �)���?4            @T@       ������������������������       �        3             T@        ������������������������       �                     �?                                 �?      �?	             0@                                `o@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        .             T@                                  L@      �?              @       ������������������������       �                     @                                �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                �`@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �t�b�       h�h)h,K ��h.��R�(KMKK��hb�B�  >��=���?a�a��?N�zv�?,�Ra���?�eY�eY�?M�4M�4�?�n�ᆫ?Hy�G�?�$I�$I�?�m۶m��?              �?�������?333333�?              �?      �?        w�qGܡ?�#�;��?�cj`?qV~B���?              �?UUUUUU�?�������?              �?�$I�$I�?۶m۶m�?              �?      �?        �q�q�?9��8���?              �?      �?        F]t�E�?/�袋.�?      �?        �B!��?�{����?              �?F]t�E�?]t�E]�?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?        f㛡���?M2/%��?�+�=�?�??j#a `�?|d�S��?7��XQ�?9��8���?�q�q�?;�;��?;�;��?      �?        �9�s��?�c�1��?��N��N�?�؉�؉�?      �?      �?              �?      �?              �?        �������?333333�?      �?      �?              �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�s�9��?�1�c��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?�������?�������?              �?�q�q�?�q�q�?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        O#,�4��?a���{�?      �?        ]t�E�?t�E]t�?      �?        �������?�������?              �?�m۶m��?�$I�$I�?333333�?�������?      �?                      �?      �?        �&M�4i�?[�lٲe�?�s�9�?c�1�c�?�A�A�?��+��+�?����?�Q�/��?����?��Ǐ?�?W�+�ɵ?�����F�?Y�B��?���7���?�{a���?GX�i���?              �?�������?�������?      �?      �?      �?                      �?              �?�?<<<<<<�?UUUUUU�?�������?�������?333333�?      �?                      �?              �?              �?      �?                      �?              �?      �?      �?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?(������?l(�����?UUUUUU�?�������?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?]t�E]�?�E]t��?              �?9��8���?�8��8��?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���Ѻ?]ʥ\ʥ�?�������?�������?�a�+�?��sK���?              �?      �?      �?�x+�R�?:�&oe�?              �?      �?        ]t�E�?t�E]t�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?      �?                      �?      �?              �?        �q�q�?r�q��?      �?        UUUUUU�?�������?              �?      �?        ?C�����?�y��`^�?T�싨��?V�	���?��VC��?�@*9/��?{�G�z�?���Q��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�-��-��?i�i��?�$I�$I�?۶m۶m�?h/�����?	�%����?              �?�?�������?�������?�������?      �?      �?              �?      �?                      �?              �?      �?      �?      �?      �?      �?                      �?      �?      �?              �?      �?        ���)k��?��)kʚ�?      �?        �o��o��?5H�4H��?'�l��&�?m��&�l�?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?      �?      �?                      �?�?�������?              �?�������?333333�?              �?      �?      �?      �?                      �?              �?X�i���?O#,�4��?�������?�������?              �?      �?        �V�9�&�?:�&oe�?�������?�������?��y��y�?�a�a�?�������?�������?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        |a���?	�=����?      �?        �N��N��?vb'vb'�?      �?      �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?��=��=�?�!�!�?���¯�?~5&��?"5�x+��?�V�9�&�?�G�z�?���Q��?*�Y7�"�?к����?      �?              �?      �?      �?        �������?UUUUUU�?              �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?-���b�?X:Ɂ���?�������?�������?      �?        ى�؉��?�؉�؉�?              �?�������?UUUUUU�?      �?        333333�?�������?              �?      �?        ��5!({�?�	A����?��^o��?��F($�??��W�?����?X�<ݚ�?�����H�?      �?                      �?      �?      �?�������?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?              �?      �?              �?      �?        �������?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJՆ�}hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@C         �                    �?SH7�j�?H           ��@              y                    �?��~а�?H           �@              6       	          pff�?84��ee�?�            pv@                      
             �?�s��:��?[             c@               
                   �_@z\�3�?-            �S@               	                    �?�g�y��?             ?@                                   �N@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     9@                                   �?�q�q��?             H@                                   �?      �?              @        ������������������������       �                     @                                  `a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                   @K@�z�G��?             D@        ������������������������       �                     ,@                                  `a@��
ц��?             :@                                  �?�d�����?             3@        ������������������������       �                      @                                   l@�eP*L��?             &@        ������������������������       �                     @                      	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               !                    �?F�����?.            @R@                                     N@�ՙ/�?             5@                                  �G@և���X�?             ,@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        "       #                   �Y@�θ�?#             J@        ������������������������       �                      @        $       '                    �H@z�G�z�?"             I@        %       &                    �?P���Q�?             4@       ������������������������       �                     3@        ������������������������       �                     �?        (       1                   @E@�z�G��?             >@        )       0       	          @33�?�eP*L��?             &@       *       +                    _@      �?             $@        ������������������������       �                     @        ,       -                    �?����X�?             @        ������������������������       �                     �?        .       /                    �N@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        2       3                    �?�S����?             3@       ������������������������       �                     *@        4       5                   �_@      �?             @        ������������������������       �                     @        ������������������������       �                     @        7       H                    �? ���g=�?�            �i@        8       ;                   @h@8^s]e�?             =@        9       :       	          `ff@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        <       A                   �`@�q�q�?             8@        =       >                    �?�q�q�?             (@        ������������������������       �                      @        ?       @       	             �?���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        B       G                    �?�8��8��?	             (@        C       F                    @O@�q�q�?             @       D       E                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        I       l                    c@��;M��?t            @f@       J       ]                   p`@H�!b	�?j            @d@       K       P                    �?������?L             [@        L       O       	             �?�C��2(�?             &@        M       N                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        Q       R                    �?`�E���?D            @X@       ������������������������       �        0            �P@        S       X       	             @��S�ۿ?             >@       T       W                   �j@ �q�q�?             8@        U       V                    X@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     *@        Y       \                    �L@r�q��?             @        Z       [                   @X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ^       c                   �`@h�WH��?             K@        _       b                   po@���Q��?             @       `       a       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        d       g       
             �?@9G��?            �H@        e       f                   @X@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        h       i                   �m@ qP��B�?            �E@       ������������������������       �                     8@        j       k                   �m@�}�+r��?
             3@        ������������������������       �                     �?        ������������������������       �        	             2@        m       n                    �F@     ��?
             0@        ������������������������       �                      @        o       p                    �?X�Cc�?             ,@        ������������������������       �                     @        q       r                    Z@�eP*L��?             &@        ������������������������       �                      @        s       v       
             �?�q�q�?             "@        t       u                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        w       x                    �J@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        z       �                    �?�m�&��?d            �b@        {       |                   Pj@�t����?-             Q@       ������������������������       �        "            �I@        }       �                   �`@��.k���?             1@        ~                          �w@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                     R@ 7���B�?7            @T@       �       �       
             �?�(\����?6             T@       ������������������������       �        .            �Q@        �       �                   �`@z�G�z�?             $@       ������������������������       �                     @        �       �                   �p@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�2Mg���?            �y@       �       �                    �?��>��?�            �t@       �       �                    �?v���a�?�            @r@        �       �                    �?���X�?&             L@        �       �                   �^@���Q��?             4@        ������������������������       �                     �?        �       �                   �e@p�ݯ��?             3@       �       �       
             �?�t����?             1@        �       �                   �e@���Q��?             @       �       �                    �?      �?             @       �       �                     L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �d@r�q��?             (@        �       �                   �m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?tk~X��?             B@        ������������������������       �                     "@        �       �                   Pb@������?             ;@        �       �                   @]@      �?             (@        ������������������������       �                     @        �       �                   �]@      �?              @        ������������������������       �                     @        �       �                    q@���Q��?             @       �       �       	          hff�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     L@��S�ۿ?             .@       ������������������������       �        	             *@        �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�n%����?�            �m@        �       �       	          ����?` A�c̭?8             Y@       ������������������������       �        ,             U@        �       �                    �?     ��?             0@       �       �                   @q@�����H�?             "@       ������������������������       �                     @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?����X�?             @       �       �                   �h@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?�����?Y             a@        �       �       	          `ff�?����X�?             <@       �       �                   �e@���|���?             6@       �       �                   �\@��.k���?             1@        ������������������������       �                     @        �       �                   �p@���!pc�?	             &@       �       �       	          ����?�����H�?             "@        �       �                    ^@      �?             @       �       �                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pt@�X�<ݺ?E             [@       �       �                   �a@��FM ò?C            @Z@        ������������������������       �                    �C@        �       �                   `p@�FVQ&�?*            �P@       �       �                   �a@�ʈD��?            �E@        ������������������������       �                     �?        �       �                   @n@@4և���?             E@       �       �                    @��?^�k�?            �A@       ������������������������       �                     A@        ������������������������       �                     �?        �       �                   �n@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     7@        �       �                   u@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `R@�p ��?            �D@        ������������������������       �                     (@        �       �                   @`@8^s]e�?             =@        ������������������������       �                     @        �       �                   �b@z�G�z�?             9@        ������������������������       �                     (@        �       �                    k@�n_Y�K�?             *@       ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @L@�w�r��?-            @S@        �       �       	             @��+��?            �B@       �       �       
             �?d��0u��?             >@       �       �                    �?     ��?             0@        ������������������������       �                      @        �       �                   �h@d}h���?
             ,@        ������������������������       �                      @        �       �                     H@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @        �       
                   @z�G�z�?             D@       �                         �`@$G$n��?            �B@       �                           R@�FVQ&�?            �@@       �             	             �?      �?             @@        �                          @`@�C��2(�?             &@       ������������������������       �                     "@                                �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     �?                    	          ����?      �?             @        ������������������������       �                      @              	                   �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 @Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  ���t��?�~�E)�?}>�����?a0��?H�k�f�?�[)J���?�k(���?��k(��?h *�3�?��jq��?�B!��?��{���?UUUUUU�?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?333333�?ffffff�?              �?�؉�؉�?�;�;�?y�5���?Cy�5��?              �?]t�E�?t�E]t�?              �?      �?      �?      �?                      �?      �?        �P�B�
�?�^�z���?�a�a�?�<��<��?�$I�$I�?۶m۶m�?              �?      �?                      �?ى�؉��?�؉�؉�?              �?�������?�������?ffffff�?�������?      �?                      �?ffffff�?333333�?]t�E�?t�E]t�?      �?      �?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?(������?^Cy�5�?      �?              �?      �?      �?                      �?ہ�v`��?��(�3J�?	�=����?|a���?�������?�������?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?Y�JV���?զ6��M�?�����H�?b�2�tk�?�q�q�?�q�q�?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?����??��W�?              �?�?�������?UUUUUU�?�������?F]t�E�?]t�E�?      �?                      �?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?B{	�%��?��^B{	�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        9/���?������?UUUUUU�?�������?      �?                      �?�}A_З?��}A�?              �?(�����?�5��P�?      �?                      �?      �?      �?      �?        �m۶m��?%I�$I��?              �?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?              �?      �?        p�j:�?�?��8��?�?<<<<<<�?              �?�?�������?�$I�$I�?۶m۶m�?              �?      �?        ffffff�?333333�?              �?      �?        h/�����?	�%����?�������?333333�?              �?�������?�������?              �?      �?      �?              �?      �?              �?        �6$oC��?��!y�?�����?��'��?ٲe˖-�?�4iҤI�?۶m۶m�?I�$I�$�?333333�?�������?              �?^Cy�5�?Cy�5��?�������?�������?�������?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?r�q��?9��8���?      �?        B{	�%��?{	�%���?      �?      �?      �?              �?      �?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�?      �?              �?      �?      �?                      �?'u_[�?�V'u�?
ףp=
�?���Q��?      �?              �?      �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?xxxxxx�?�$I�$I�?�m۶m��?F]t�E�?]t�E]�?�?�������?              �?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?      �?      �?      �?      �?                      �?      �?              �?                      �?              �?              �?��8��8�?�q�q�?��~���?8�8��?      �?        >����?|���?A_���?�}A_з?              �?n۶m۶�?�$I�$I�?_�_��?�A�A�?      �?                      �?�m۶m��?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        8��18�?dp>�c�?              �?|a���?	�=����?              �?�������?�������?      �?        ;�;��?ى�؉��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?
qV~B��?{����1�?�S�n�?*�Y7�"�?DDDDDD�?wwwwww�?      �?      �?      �?        ۶m۶m�?I�$I�$�?              �?      �?      �?      �?                      �?      �?                      �?ffffff�?ffffff�?���L�?к����?|���?>����?      �?      �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�$"hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�@         d       	          ����?�>�Ļ`�?I           ��@               /       
             �?@jn�lo�?           `{@               .                   �a@DS���|�?[             a@                                  �?�`�=	�?F            �Y@               
                     G@�n_Y�K�?             *@               	       	          ����?�q�q�?             @                                 �[@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                  �d@؇���X�?             @                                   `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               '                   �`@ףp=
�?>            �V@              "                   xr@P���Q�?8             T@                     	          833�?P�Lt�<�?5             S@                                 @W@ ��PUp�?1            �Q@                                 �^@�(\����?             D@                                 `]@ ��WV�?             :@        ������������������������       �                     *@                                   �?$�q-�?
             *@       ������������������������       �                     $@                                   �?�q�q�?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     ?@                !                   (p@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        #       &                    �?      �?             @       $       %                   �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        (       -                    �?      �?             $@       )       ,                     @����X�?             @       *       +                    X@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     A@        0       C                    �K@�iD���?�            �r@       1       2       	          ���ٿ�IєX�?�            �k@        ������������������������       �                     �?        3       B                    �?�1�`jg�?�            �k@        4       9                    �?V�a�� �?"             M@        5       6                   �i@      �?             ,@        ������������������������       �                     @        7       8                     D@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        :       ;                    X@�Ra����?             F@        ������������������������       �                      @        <       =                    �I@@4և���?             E@       ������������������������       �                     B@        >       A                    @J@      �?             @       ?       @                   0c@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        i            @d@        D       c                   xt@H�z���?3             T@       E       N                   �T@N��c��?1            @S@        F       M                   �c@�q�q�?             (@       G       L                    �?����X�?             @        H       I                    �?�q�q�?             @        ������������������������       �                     �?        J       K                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        O       Z       	          ����?�z����?)            @P@       P       W                   �r@8��8���?             H@       Q       V                    �?��Y��]�?            �D@        R       S                   `b@$�q-�?             *@       ������������������������       �                     &@        T       U                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     <@        X       Y                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        [       `                    �?ҳ�wY;�?             1@        \       ]                   Ph@�q�q�?             @        ������������������������       �                     �?        ^       _                    �P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        a       b                    �M@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        e       �                    �?�G�z.�?/            ~@       f       �                   0e@�-�j���?�             t@       g       �                   �u@l{��b��?�            �s@       h       w                   @\@��GEI_�?�            s@        i       j                   @Y@>A�F<�?             C@        ������������������������       �        	             (@        k       v       
             �?R�}e�.�?             :@       l       q                     M@b�2�tk�?             2@       m       n                   �]@���Q��?             $@        ������������������������       �                     @        o       p       	          033@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        r       s                   �^@      �?              @        ������������������������       �                     @        t       u                   @h@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        x       �                    �R@�7,��?�            �p@       y       z                    @H@�w�>τ�?�            pp@        ������������������������       �                     E@        {       �                    �?��s97�?�            �k@        |       }                   �c@     ��?#             P@       ������������������������       �                     I@        ~              
             �?@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        �       �                    �?�B�ǈ�?g            �c@       �       �                    c@,���$�?@            @X@       �       �                    �? p�/��?:            @V@        �       �                   xr@�r����?	             .@       ������������������������       �                     *@        ������������������������       �                      @        �       �                    �?�?�|�?1            �R@        �       �                   0n@z�G�z�?             @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   p`@@	tbA@�?-            @Q@       ������������������������       �        #             I@        �       �       
             �?�}�+r��?
             3@       ������������������������       �                     *@        �       �                   Pa@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                    @N@      �?             @        ������������������������       �                      @        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?P���Q�?'             N@        �       �       
             �?8�Z$���?	             *@        �       �                    @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?�C��2(�?             &@       �       �                   @_@�����H�?             "@       ������������������������       �                     @        �       �                    �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?`Ql�R�?            �G@        �       �                    �L@      �?              @        �       �                   �^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �C@        �       �       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?���|���?             &@       �       �                    b@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �H@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�j����?g            �c@       �       �                   �b@��Cp]�?F            �\@        �       �                    �?��WV��?             J@        �       �                   �b@�����H�?
             2@       ������������������������       �                     .@        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     P@h+�v:�?             A@       �       �                   Pb@�q�����?             9@       �       �                   0b@�ՙ/�?             5@       �       �                   @g@��S���?	             .@       �       �                    \@      �?              @        ������������������������       �                     @        �       �       	          @33�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?����X�?+            �O@        ������������������������       �                     5@        �       �                   ``@և���X�?             E@       �       �                    �?      �?             8@       �       �                    @F@      �?             0@        �       �                   Pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    m@      �?              @       ������������������������       �                     @        �       �                   �^@      �?             @       �       �                   @p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �L@�q�q�?             2@        �       �                   m@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �n@r�q��?             (@       �       �                   �a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �c@�%^�?!            �E@        ������������������������       �                     (@        �       �                    �J@f���M�?             ?@        �       �                   c@r�q��?             @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    Y@�+e�X�?             9@        ������������������������       �                     �?        �       �       	          ����?�q�q�?             8@        �       �                    �P@      �?              @       �       �                   8v@�q�q�?             @       �       �                    �L@z�G�z�?             @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �                           @      �?             0@       ������������������������       �        	             *@                                �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B0  Qm4��?X��;�?zH�!���?o3����?�uy)�?I�ܺ�?�H%�e�?��6���?ى�؉��?;�;��?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?              �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?�������?�������?�������?ffffff�?(�����?���k(�?��V،?��ۥ���?�������?333333�?;�;��?O��N���?              �?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?              �?              �?�������?�������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?�������?UUUUUU�?              �?      �?                      �?              �?              �?Of�b�?;��ϼ�?�?�?              �?A��)A�?�־a�?��{a�?a���{�?      �?      �?              �?      �?      �?              �?      �?        ]t�E]�?]t�E�?              �?n۶m۶�?�$I�$I�?      �?              �?      �?�������?333333�?      �?                      �?      �?              �?        �������?�������?�����?5�wL��?�������?�������?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?[��Z���?�Z��Z��?�������?�������?8��18�?������?�؉�؉�?;�;��?      �?              �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        /�袋.�?F]t�E�?              �?      �?                      �?ffffff�?ffffff�?(�ˀO�?��6�?�&��jq�?${�ґ�?;ڼOqɰ?�d����?Cy�5��?������?              �?�;�;�?'vb'vb�?9��8���?�8��8��?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�!�c��?��y#q�?\�Nj�?�~k^��?              �?�{�{�?�@h�@h�?      �?     ��?              �?�$I�$I�?n۶m۶�?              �?      �?        �n�{DN�?$r�p7��?���fy�?�,O"Ӱ�?p�\��?�G?�я�?�?�������?              �?      �?        к����?*�Y7�"�?�������?�������?      �?      �?      �?                      �?              �?ہ�v`��?�%~F��?              �?(�����?�5��P�?              �?UUUUUU�?�������?      �?                      �?      �?      �?              �?333333�?�������?      �?      �?      �?              �?      �?      �?                      �?              �?�������?ffffff�?;�;��?;�;��?      �?      �?              �?      �?        F]t�E�?]t�E�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?              �?W�+�ɕ?}g���Q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?      �?                      �?F]t�E�?]t�E]�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?UUUUUU�?      �?                      �?n���7�?${�ґ�?I�ø_��?m5x�@��?��؉���?��N��N�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        xxxxxx�?�������?�p=
ף�?���Q��?�<��<��?�a�a�?�������?�?      �?      �?      �?              �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?              �?�m۶m��?�$I�$I�?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?      �?      �?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?�������?333333�?              �?      �?                      �?�}A_�?�}A_��?              �?��Zk���?��RJ)��?�������?UUUUUU�?      �?      �?      �?                      �?      �?        ���Q��?R���Q�?      �?        �������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?              �?                      �?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJK55EhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKۅ�h��B�6         �       
             �?������?6           ��@              #                    �F@�H"ȏ��?4           @                                   �?�A����?1            �T@                                  �?h�WH��?              K@                                   `@      �?              @        ������������������������       �                      @               
                    �?r�q��?             @              	                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                  pb@�nkK�?             G@                                  �?�Ń��̧?             E@                                  pb@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     B@                                   �C@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                      	          ����?X�Cc�?             <@                                  `a@      �?             0@                                  @`@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                   m@�<ݚ�?             "@                                  �f@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                   �o@r�q��?
             (@       ������������������������       �                     "@        !       "                   �d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        $       /       	          ����?ЖkÄ�?           �y@        %       (       
             �?@3����?>             [@        &       '                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        )       *                   �p@�ջ����?;             Z@       ������������������������       �        4            �V@        +       .                    �?$�q-�?             *@        ,       -                   (r@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        0       a                    �?�=��=��?�            0s@       1       V                   �a@4�f����?�             l@       2       I                   pr@ �	.��?X            ``@       3       6       	          ����?@-�_ .�?K            �[@        4       5                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        7       F                    c@ '��h�?I            @[@       8       E                    �L@`�(c�?B            �X@       9       :       	          ����? �h�7W�?#            �J@        ������������������������       �                     �?        ;       @                   @X@ ��WV�?"             J@        <       =                   �Y@�q�q�?             @        ������������������������       �                     �?        >       ?                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        A       D                    �?@�E�x�?            �H@        B       C                   h@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     F@        ������������������������       �                    �F@        G       H                   `c@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        J       O                    s@��Q��?             4@        K       N       	             �?����X�?             @       L       M                   �r@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        P       Q       	          ����?8�Z$���?	             *@        ������������������������       �                     �?        R       S                   `v@�8��8��?             (@       ������������������������       �                     "@        T       U                   �x@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        W       \                   �r@��V�I��?5            �W@       X       [                    �?��'�`�?.            �T@        Y       Z                   pl@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        )            �S@        ]       ^                   �c@"pc�
�?             &@        ������������������������       �                     @        _       `                   �s@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        b       g                    �?yÏP�?8            �T@        c       f       	          ����?      �?             0@        d       e                    Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        h       k       
             �?�X����?-            �P@        i       j                   �]@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        l       w       	             �?^(��I�?&            �K@        m       n                   Pk@��S���?             .@        ������������������������       �                     @        o       v                    �?�z�G��?             $@       p       u                    o@���Q��?             @       q       r                   �a@�q�q�?             @        ������������������������       �                     �?        s       t                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        x       �       	          ���@z�G�z�?             D@       y       z                   �Q@     ��?             @@        ������������������������       �                     @        {       |                   �[@\-��p�?             =@        ������������������������       �                      @        }       �                    @J@�>����?             ;@        ~                          c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���N8�?             5@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             2@        ������������������������       �                      @        �       �                    �?H���0��?           Pz@       �       �                   �O@�ˠTX�?�             v@        �       �                    �?�z�G��?             4@       �       �       	          ����?���Q��?
             $@       �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    @L@��{�J �?�            �t@       �       �                    �I@XB���?�            Pp@       �       �                    �? ������?r            �g@        �       �                   @^@�˹�m��?             C@        �       �       	          ����?z�G�z�?	             .@       �       �                   �q@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        ������������������������       �        Z            �b@        �       �                   �g@�8��8��?,             R@       �       �                   �d@�nkK�?+            @Q@       ������������������������       �        #             K@        �       �                   �_@z�G�z�?             .@        �       �                    �J@և���X�?             @        �       �                   �p@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �M@�ګH9�?*            �Q@        �       �                    �?��>4և�?             <@       �       �                   `b@�G��l��?             5@       �       �                    �?d}h���?
             ,@        �       �                   �d@���Q��?             @        ������������������������       �                      @        �       �                   0f@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@�����H�?             "@        �       �                    @M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `c@�T|n�q�?            �E@       ������������������������       �                     :@        �       �                    �?j���� �?
             1@       �       �                    �?r�q��?             (@        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?�q�q�?)            @Q@       �       �       	          ����?      �?"             N@        �       �                   Pd@X�<ݚ�?             ;@       �       �                   0a@�LQ�1	�?             7@       �       �                    @N@�t����?	             1@       ������������������������       �                     $@        �       �                   �o@����X�?             @        ������������������������       �                     @        �       �                    @Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    c@�C��2(�?            �@@       �       �                    S@h�����?             <@        �       �       	          `ff�?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     8@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          033�?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �#@y��?'�_|C��?얋͒�?E��L�?�18���?�cp>�?B{	�%��?��^B{	�?      �?      �?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?d!Y�B�?�Mozӛ�?�a�a�?��<��<�?UUUUUU�?�������?              �?      �?                      �?      �?      �?              �?      �?        %I�$I��?�m۶m��?      �?      �?۶m۶m�?�$I�$I�?              �?      �?        �q�q�?9��8���?�������?333333�?              �?      �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        :�3�X�?r�����?h/�����?���Kh�?      �?      �?      �?                      �?;�;��?;�;��?              �?;�;��?�؉�؉�?�������?�������?      �?                      �?              �?P�A�C�?��/��?߼�xV4�?d��0u��?�U���g�?@u���?к����?S�n0E�?      �?      �?      �?                      �?�w� z|�?���]8��?և���X�?��)x9�?"5�x+��?��sHM0�?      �?        ;�;��?O��N���?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        9/���?և���X�?�������?�������?      �?                      �?              �?              �?F]t�E�?/�袋.�?      �?                      �?ffffff�?�������?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?AL� &W�?<�����?��k���?1P�M��?�������?�������?      �?                      �?              �?F]t�E�?/�袋.�?              �?�������?333333�?      �?                      �?Q��+Q�?W�v%jW�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ]t�E]�?�E]t��?]t�E]�?F]t�E�?              �?      �?        J��yJ�?�7�}���?�������?�?              �?ffffff�?333333�?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        ffffff�?ffffff�?      �?      �?      �?        �{a���?a����?      �?        h/�����?�Kh/��?UUUUUU�?�������?              �?      �?        �a�a�?��y��y�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?<���c�?�-шs�?F]t�E�?�E]tѽ?333333�?ffffff�?333333�?�������?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?M�_{�e�?�%�Ѵ?GX�i���?�{a���?��}��}�?AA�?��P^Cy�?^Cy�5�?�������?�������?�؉�؉�?;�;��?      �?                      �?              �?      �?              �?        UUUUUU�?UUUUUU�?�Mozӛ�?d!Y�B�?      �?        �������?�������?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?              �?              �?                      �?e�v�'��?6��9�?۶m۶m�?I�$I�$�?1�0��?��y��y�?I�$I�$�?۶m۶m�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?      �?      �?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?        ���)k��?6eMYS��?      �?        �������?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?      �?�q�q�?r�q��?d!Y�B�?Nozӛ��?�?<<<<<<�?              �?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?      �?              �?        F]t�E�?]t�E�?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?�������?333333�?              �?      �?        �q�q�?�q�q�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ&hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hK�)      hyMhzh)h,K ��h.��R�(KM��h��B@F         �                    �?>���i��??           ��@              I                    �?����?`           X�@                      
             �?l?Z��i�?�            `j@                     	          833�?�����?K            �[@        ������������������������       �                     E@               	       	          ����?�q�q�?/            @Q@                                   �?$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        
                          �`@����>4�?(             L@                                  hq@     ��?             @@                                 �^@ףp=
�?             4@                                  Pn@�<ݚ�?             "@                                 @[@      �?              @        ������������������������       �                     @                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@                      	          ���@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @                                  �x@ �q�q�?             8@       ������������������������       �                     4@                                   b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               "                    T@؁sF���?=             Y@               !                    �?ףp=
�?             4@                                   �\@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     0@        #       @                    �M@���Q8�?/             T@       $       9       	          ����?     8�?&             P@       %       4                    @F@�C��2(�?!            �K@        &       3                   �b@���y4F�?             3@       '       0                   �e@�t����?             1@       (       )                    �E@@4և���?	             ,@       ������������������������       �                      @        *       +                    �?r�q��?             @        ������������������������       �                      @        ,       -                   0o@      �?             @        ������������������������       �                      @        .       /                   �u@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        5       6                   �r@������?             B@       ������������������������       �                     ?@        7       8                   �d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        :       ?                    o@�q�q�?             "@       ;       >                   0e@      �?             @        <       =                   0l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        A       H       	          `ff�?      �?	             0@       B       G       	            �?z�G�z�?             .@       C       D                   �b@�q�q�?             "@        ������������������������       �                      @        E       F                   �_@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        J       �                   �g@JgƟn��?�            �u@       K       l                    �K@�k�'7��?�            `u@       L       U                   d@8���@�?�            `m@        M       R                   �`@���!pc�?             6@       N       Q                   �P@      �?             0@        O       P       	          ����?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        S       T                    @G@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        V       k       
             �?��$xtW�?�            �j@        W       b                   Pp@d,���O�?            �I@       X       Y       	            �?�#-���?            �A@        ������������������������       �                     *@        Z       a                   0m@��2(&�?             6@        [       `                   �`@      �?              @       \       _                   �\@r�q��?             @        ]       ^       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        c       d                    �?      �?	             0@        ������������������������       �                     @        e       j                   �b@r�q��?             (@       f       i                    @�C��2(�?             &@       g       h                   `\@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        k            @d@        m       �       	             @r���@�?F            �Z@       n       o       	          ���修Y �K�?>            @X@        ������������������������       �                     @        p       �                   �d@����X�?<            �V@       q       �                    �?�w�r��?4            @S@        r       }       
             �?z�G�z�?             9@        s       t       	             �?X�<ݚ�?             "@        ������������������������       �                      @        u       |                     P@և���X�?             @       v       {                   �b@�q�q�?             @       w       x                   �[@z�G�z�?             @        ������������������������       �                      @        y       z                   0m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ~                          �c@      �?
             0@       ������������������������       �                     &@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�E��
��?$             J@        �       �                    p@8����?             7@       �       �                    �L@�8��8��?             (@        �       �       
             �?z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?�eP*L��?             &@        �       �                   p`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	             �?z�G�z�?             @        ������������������������       �                      @        �       �       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          pff�?l��[B��?             =@       �       �                    \@��Q��?             4@        ������������������������       �                     �?        �       �                   pa@�����?             3@        �       �                    �M@      �?              @        �       �                   �g@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�eP*L��?             &@        �       �                    �N@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?             @       �       �                    �O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �_@      �?              @        ������������������������       �                     �?        �       �       
             �?؇���X�?             @        ������������������������       �                     @        �       �                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        �       �                    �M@ףp=
�?             $@        �       �                   `c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �i@<�,@���?�            �v@        �       �                   �b@`2U0*��?N            @_@       �       �                   �c@@3����?C             [@       �       �                   �`@@䯦s#�?A            �Z@       ������������������������       �        1             T@        �       �                    @M@ ��WV�?             :@       ������������������������       �        
             0@        �       �                   �^@ףp=
�?             $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @U@@�0�!��?             1@       �       �       
             �?�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �       	          033�?@�0�!��?�            �m@        �       �                   �n@�~8�e�?            �I@        �       �                   �k@�E��ӭ�?             2@        �       �                    �J@և���X�?             @        ������������������������       �                      @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   n@�C��2(�?             &@       ������������������������       �                     @        �       �                   @n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �r@���!pc�?            �@@       �       �                    �N@      �?             8@       �       �                    �?���7�?             6@       ������������������������       �        	             3@        �       �                     H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?Ԧ\�s�?t            `g@        �       �                    �?������?             A@       �       �                    �M@�LQ�1	�?             7@       �       �                    @H@��S�ۿ?
             .@        �       �                    �?؇���X�?             @        �       �                    @D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @b@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   po@�eP*L��?             &@        ������������������������       �                     @        �       �                   `]@؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �                          �J@�:�]��?_             c@        �                          @J@j�q����?             I@       �              	          ����?��p\�?            �D@        �       �                   �\@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                �b@�?�|�?            �B@       ������������������������       �                     >@                                 o@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                    	             @�q�q�?             "@                   	             �?���Q��?             @        ������������������������       �                     �?        	      
                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                �j@ f^8���?A            �Y@                                @_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 c@@�E�x�?<            �X@                                �R@�L��ȕ?8            @W@       ������������������������       �        6            �V@                                �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 q@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  �Q��Q��?W�W��?�Oyk���?g`)u�?Tyt�=��?V��a��?\�9	ą�?镱��^�?              �?UUUUUU�?UUUUUU�?�؉�؉�?;�;��?      �?                      �?I�$I�$�?n۶m۶�?      �?      �?�������?�������?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?�z�G��?=
ףp=�?�������?�������?      �?      �?      �?                      �?              �?�������?ffffff�?     ��?      �?]t�E�?F]t�E�?6��P^C�?(������?<<<<<<�?�?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?      �?              �?      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�q�q�?�q�q�?      �?        �������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?              �?                      �?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?                      �?              �?      �?        ��#�;�?�qG��?-����b�?Lg1��t�?�"��i�? ��§��?F]t�E�?t�E]t�?      �?      �?9��8���?�q�q�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?����?��n�?�?�������?PPPPPP�?�A�A�?_�_�?      �?        ��.���?t�E]t�?      �?      �?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?              �?      �?      �?        UUUUUU�?�������?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?      �?              �?        Ei|d��?u-7���?���
|q�?����?              �?�m۶m��?�$I�$I�?{����1�?
qV~B��?�������?�������?r�q��?�q�q�?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?        �������?�������?      �?                      �?;�;��?��؉���?d!Y�B�?8��Moz�?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ]t�E�?t�E]t�?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ���=��?GX�i���?�������?ffffff�?              �?Q^Cy��?^Cy�5�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        t�E]t�?]t�E�?�m۶m��?�$I�$I�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?9��8���?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?My�N���?��@�S��?{�G�z�?���Q��?h/�����?���Kh�?�x+�R�?R����?              �?;�;��?O��N���?              �?�������?�������?      �?      �?      �?                      �?              �?      �?      �?      �?                      �?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?ZZZZZZ�?�������?222222�?�q�q�?r�q��?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?      �?              �?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?        t�E]t�?F]t�E�?      �?      �?F]t�E�?�.�袋�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?a�2a�?�|�ٓ�?�?xxxxxx�?Y�B��?��Moz��?�?�������?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?      �?      �?              �?      �?        ]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�?}}}}}}�?
ףp=
�?=
ףp=�?��+Q��?�]�ڕ��?      �?      �?      �?                      �?к����?*�Y7�"�?              �?�$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?�������?333333�?              �?      �?      �?      �?                      �?      �?        ��VCӝ?H%�e�?�������?�������?      �?                      �?9/���?և���X�?X`��?��~���?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJd+�3hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�A         ~       	          `ff�?��J�0�?I           ��@              1       
             �?uvI��?<           �~@                                  �h@b�����?m             e@                                   �? ��WV�?1            �S@       ������������������������       �        !            �J@                                   �?H%u��?             9@                                   �H@�q�q�?             @        ������������������������       �                     �?        	       
                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?���7�?             6@                                  @M@$�q-�?             *@                                  �S@z�G�z�?             @                                  �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@               $                    �?����?<            �V@                      
             �?���>4��?             <@        ������������������������       �                     @                                   �?      �?             8@        ������������������������       �                     @               #                    �?      �?             4@                                 @^@�eP*L��?	             &@        ������������������������       �                     @                                  �c@      �?              @       ������������������������       �                     @                       	          833�?�q�q�?             @        ������������������������       �                     �?        !       "                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        %       *                    �F@��s����?'            �O@        &       '                    �?��
ц��?             *@        ������������������������       �                     @        (       )                   0o@      �?              @       ������������������������       �                     @        ������������������������       �                      @        +       0                   �e@H%u��?             I@       ,       -       	          hff�? i���t�?            �H@       ������������������������       �                    �E@        .       /                    @J@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        2       ]                    �?���G�?�            t@        3       H                    `@����?9            @V@        4       C                    �?�>$�*��?            �D@       5       >                   `]@      �?             @@       6       ;                   �b@�ՙ/�?             5@       7       :       	          433�?���Q��?             $@       8       9                   `\@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        <       =                   �f@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ?       @                    V@���!pc�?	             &@        ������������������������       �                      @        A       B                   0e@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        D       E                   �q@�<ݚ�?             "@       ������������������������       �                     @        F       G                   �r@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        I       N                    �L@r�q��?             H@       J       K                   �b@г�wY;�?             A@       ������������������������       �                     >@        L       M                   �b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        O       P                    �?      �?
             ,@        ������������������������       �                      @        Q       X                   `a@�q�q�?	             (@        R       W                    �?�q�q�?             @       S       V                   a@z�G�z�?             @       T       U                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        Y       Z                   �b@r�q��?             @       ������������������������       �                     @        [       \                    [@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ^       }                   h@�a�� �?�             m@       _       r                    @x���a�?�            �l@       `       q                   �c@�J�T�?�            �j@       a       h                   �b@����˵�?M            �]@       b       g                   �_@��F�D�?>            �X@        c       f                   @c@�8��8��?             8@        d       e                   @^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        ������������������������       �        -            �R@        i       l                    �?���y4F�?             3@       j       k                    �?�r����?             .@        ������������������������       �                      @        ������������������������       �        
             *@        m       n       	          �����      �?             @        ������������������������       �                     �?        o       p                   @Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        @            �W@        s       |                    �M@      �?             0@       t       u                    h@և���X�?             @        ������������������������       �                     �?        v       w                   �j@�q�q�?             @        ������������������������       �                     @        x       {       	          ����?�q�q�?             @       y       z                    o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @               �                   �c@�7�ɣ�?           �z@       �       �                    �?��X@�?�            �v@       �       �                   �m@��S�ۿ?�            �p@       �       �                    �?Pt�nٔ�?l            �e@       �       �                    c@ d�=��?D            @\@       �       �                   �Z@      �?C             \@        �       �                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�1�`jg�?A            �[@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                     M@      �?             @        ������������������������       �                      @        �       �                   �R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��9J���?<             Z@       �       �                     E@ ��N8�?/             U@        �       �       	          ����?�8��8��?             (@        ������������������������       �                      @        �       �                    @D@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        *             R@        �       �                    @L@ףp=
�?             4@        ������������������������       �                     "@        �       �       	          ����?"pc�
�?             &@        �       �                    �O@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        (             N@        �       �                   0c@�^'�ë�?@            @X@       �       �                    �J@     ��??             X@        �       �                    �?�MI8d�?            �B@        �       �                   �^@���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?     ��?             @@       ������������������������       �                     8@        �       �                    �?      �?              @       �       �                     H@      �?             @        ������������������������       �                      @        �       �                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   @Z@����˵�?)            �M@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �       	          033�? �Jj�G�?&            �K@        ������������������������       �                     6@        �       �                    �?Pa�	�?            �@@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        ������������������������       �                     �?        �       �                   �n@$�ݏ^��?7            �V@       �       �                    `@:2vz�M�?%            �N@       �       �                   0j@������?             A@       �       �                    �P@���N8�?             5@       ������������������������       �        
             .@        �       �       	          hff@r�q��?             @       �       �                   �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �Q@��
ц��?             *@       �       �                   P`@�z�G��?             $@        ������������������������       �                     @        �       �                   �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @N@�q�q�?             ;@       �       �       	             @      �?             2@       �       �                    �?�	j*D�?
             *@        ������������������������       �                     @        �       �                    �?և���X�?             @       �       �                    �?���Q��?             @       �       �                   �a@�q�q�?             @        ������������������������       �                     �?        �       �                     H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   �b@ܷ��?��?             =@       �       �                   @^@ 7���B�?             ;@        �       �       	          ����?؇���X�?             @        �       �                   `c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                      @        �       �                    �?      �?*             Q@       �       �                    �L@x�K��?!            �I@       �       �                    `@      �?             B@       �       �       	          ���@�G�z��?             4@       �       �       	          ����?������?             .@        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                     E@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �        
             0@        �       �                    �?������?	             .@       �       �                    �?ףp=
�?             $@        �       �                   �c@      �?             @       �       �       	          `ff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �_@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                          pi@@�0�!��?	             1@        ������������������������       �                      @                    	             @��S�ۿ?             .@                                �?      �?              @                                �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��hb�Bp  �̓"��?�6�n��?��X��?
^N��)�?g\�5�?@�(ݾ��?;�;��?O��N���?              �?���Q��?)\���(�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        F]t�E�?�.�袋�?;�;��?�؉�؉�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?R�Q��?Ws5Ws5�?n۶m۶�?I�$I�$�?      �?              �?      �?      �?              �?      �?]t�E�?t�E]t�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�a�a�?z��y���?�؉�؉�?�;�;�?              �?      �?      �?      �?                      �?���Q��?)\���(�?����X�?/�����?              �?�������?UUUUUU�?              �?      �?              �?        �v����?�$RY���?NmjS���?e%+Y�J�?�����?�18���?      �?      �?�a�a�?�<��<��?333333�?�������?۶m۶m�?�$I�$I�?      �?                      �?              �?F]t�E�?/�袋.�?              �?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?                      �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?�?�?      �?              �?      �?      �?                      �?      �?      �?      �?        �������?�������?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        sO#,�4�?��=���?�_OE��?��
�[�?(�K=�?��V؜?W'u_�?��/���?j�J�Z�?[�R�֯�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        6��P^C�?(������?�������?�?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?2�ީk9�?�_����?a�`��?(}�'}��?�?�������?���"��?4�q�-��?x�!���?���	��?      �?      �?      �?      �?              �?      �?        �־a�?A��)A�?      �?      �?              �?      �?      �?      �?              �?      �?              �?      �?        �؉�؉�?;�;��?�a�a�?�y��y��?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?�������?�������?              �?F]t�E�?/�袋.�?      �?      �?      �?                      �?              �?      �?                      �?���Id�?=�L�v��?      �?      �?L�Ϻ��?��L���?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?      �?      �?      �?      �?      �?              �?      �?      �?                      �?              �?��/���?W'u_�?      �?      �?      �?                      �?��)A��?k߰�k�?              �?|���?|���?      �?      �?      �?                      �?              �?      �?        �I��I��?[�[��?��!XG�?��6�S\�?�?xxxxxx�?�a�a�?��y��y�?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�;�;�?�؉�؉�?ffffff�?333333�?      �?              �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?vb'vb'�?;�;��?      �?        ۶m۶m�?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?              �?      �?        a���{�?��=���?h/�����?	�%����?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?              �?      �?ssssss�?�?      �?      �?�������?�������?wwwwww�?�?�������?333333�?              �?      �?        �������?�������?              �?      �?                      �?      �?        �?wwwwww�?�������?�������?      �?      �?      �?      �?      �?                      �?              �?              �?333333�?�������?              �?      �?        �������?ZZZZZZ�?      �?        �?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���2hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�B         �       	          033�?~jÚʞ�?J           ��@                                 `^@^�K����?=            @                      
             �?�	j*D�?H             Z@                                 �W@l��\��?,             Q@        ������������������������       �                     5@                                  m@��E�B��?            �G@                                  �L@�MI8d�?            �B@                                 0l@����X�?             5@       	                          �`@���y4F�?             3@       
              	          033�?�	j*D�?             *@                                 �X@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     $@                      	          ����?�E��ӭ�?             B@                                  @O@؇���X�?             <@                     	             �`2U0*��?             9@        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?                      	          hff�?؇���X�?             @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                K                    �?BTӓ�=�?�            �x@        !       "                   �_@�����'�?I            @]@        ������������������������       �                     9@        #       4                    �?��*(��?:             W@        $       3       	          ����?     ��?             @@       %       ,                   �p@�n_Y�K�?             :@       &       '                   �i@�q�q�?             (@        ������������������������       �                      @        (       )                    �?z�G�z�?             $@       ������������������������       �                     @        *       +       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        -       2                    �O@؇���X�?             ,@       .       1                    �L@$�q-�?             *@        /       0                    �I@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        5       J       	          ����?��Q��?(             N@       6       ;                    �?(옄��?             G@        7       8                   �b@      �?              @        ������������������������       �                     @        9       :       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        <       =                   0e@D�n�3�?             C@        ������������������������       �                     @        >       I                   �a@�'�=z��?            �@@       ?       @                   �f@`�Q��?             9@        ������������������������       �                      @        A       F                     D@��+7��?             7@        B       C                    @A@�q�q�?             @        ������������������������       �                     �?        D       E                   @_@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        G       H       
             �?�t����?             1@        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                      @        ������������������������       �        
             ,@        L       g                    @L@p��R(�?�            Pq@       M       N                    I@��qn�H�?�            �i@        ������������������������       �                     @        O       f                   @g@���a�\�?�            @i@       P       W                   Pn@�X�� �?�             i@       Q       V                   `c@�Ru߬Α?K            �\@        R       U                    �?      �?             @        S       T                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        G            �[@        X       a       
             �?�ʈD��?7            �U@        Y       `                    �?և���X�?             ,@       Z       [                    �?���!pc�?             &@        ������������������������       �                     @        \       _                    �?���Q��?             @       ]       ^                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        b       e                   0c@������?/             R@        c       d                   �n@�����H�?             2@        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �        #             K@        ������������������������       �                      @        h       {                    @v���EO�?&            �Q@       i       j                    �?V�a�� �?             M@        ������������������������       �                     1@        k       v       	            �?������?            �D@       l       q                   Pc@z�G�z�?             >@       m       p                    @M@�KM�]�?
             3@        n       o       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     .@        r       u                    c@���|���?             &@       s       t                    �N@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        w       x                    �L@�eP*L��?             &@        ������������������������       �                     @        y       z                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        |       }                   �a@�n_Y�K�?             *@        ������������������������       �                     @        ~       �                    �?r�q��?             @               �                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �b@����K�?           @z@       �       �                   P`@�-q���?�            �u@        �       �                   @r@�n`���?d            `c@       �       �                   �^@���V��?V            �`@        �       �                   �X@ ,��-�?%            �M@        �       �                    @P@8�Z$���?             *@       �       �                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�nkK�?             G@        ������������������������       �                     �?        �       �                    �?����?�?            �F@       ������������������������       �                    �A@        �       �                    @K@ףp=
�?             $@        �       �       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�A+K&:�?1             S@       �       �                   �_@�����H�?"             K@        �       �       	             �?�q�q�?             @        ������������������������       �                      @        �       �                   �k@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �F@�8��8��?             H@        ������������������������       �                     0@        �       �       	          ����?      �?             @@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?@4և���?             <@       �       �                     K@�nkK�?             7@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �       �                    ]@z�G�z�?             @        ������������������������       �                      @        �       �                   @_@�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �m@      �?             6@       �       �                   `U@�θ�?
             *@        ������������������������       �                      @        �       �                    �?�C��2(�?             &@        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �       	          ����?r�q��?             @        ������������������������       �                     @        �       �                   @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @_@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�G�z��?             4@       �       �       	          `ff�?���Q��?             .@       �       �                   @X@      �?             (@        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                    �K@����X�?             @       �       �                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?p�qG�?z             h@        �       �                    �?�<ݚ�?             2@       �       �       	             �?@4և���?	             ,@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   po@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        �       �                    \@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pv@XB���?m            �e@       �       �                   �h@�Sa��?i            �d@        �       �                   �e@�1�`jg�?!            �K@       �       �                   �c@�O4R���?             �J@       ������������������������       �                     C@        �       �       
             �?��S�ۿ?	             .@       ������������������������       �                     (@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        H             \@        �       �       
             �?և���X�?             @       �       �                    a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �L@�Jhu4��?/            @R@       �       �                   �c@�GN�z�?             F@        �       �                   `j@��S���?             .@        ������������������������       �                     @        �       �                    �G@�q�q�?             (@        �       �                   c@�q�q�?             @        �       �                   �u@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   `a@ܷ��?��?             =@       �       �       	          ����?���7�?             6@        ������������������������       �                     �?        ������������������������       �                     5@        �       �                   �e@����X�?             @        ������������������������       �                     @        �       �       	          pff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    c@8^s]e�?             =@        ������������������������       �                     @        �       
                  xu@z�G�z�?             9@                                 �?r�q��?             8@       ������������������������       �                     .@              	      	          `ff@X�<ݚ�?             "@                               �q@����X�?             @                                �?r�q��?             @                                b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  g�����?L��/��?��q���?����?;�;��?vb'vb'�?�������?------�?              �?AL� &W�?�l�w6��?L�Ϻ��?��L���?�$I�$I�?�m۶m��?(������?6��P^C�?;�;��?vb'vb'�?      �?      �?      �?                      �?      �?                      �?      �?                      �?              �?�q�q�?r�q��?۶m۶m�?�$I�$I�?���Q��?{�G�z�?              �?      �?                      �?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?yG5����?q�)`>�?۬�ڬ��?�)��)��?              �?��,d!�?���7���?      �?      �?ى�؉��?;�;��?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?;�;��?�؉�؉�?�������?�������?              �?      �?                      �?      �?                      �?�������?ffffff�?���,d�?ӛ���7�?      �?      �?              �?      �?      �?              �?      �?        l(�����?(������?      �?        |��|�?|���?��(\���?{�G�z�?              �?zӛ����?Y�B��?UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?        <<<<<<�?�?              �?      �?                      �?      �?        0���M�?�#�?24��~��?r^�	��?              �?D�I��A�?��g���?���(\��?
ףp=
�?���#��?p�}��?      �?      �?      �?      �?              �?      �?              �?              �?        A_���?�}A_з?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�q�q�?�q�q�?�q�q�?�q�q�?              �?      �?              �?                      �?�
��V�?�ԓ�ۥ�?��{a�?a���{�?      �?        �v%jW��?��+Q��?�������?�������?�k(���?(�����?      �?      �?              �?      �?              �?        ]t�E]�?F]t�E�?9��8���?�q�q�?      �?                      �?              �?]t�E�?t�E]t�?              �?�������?UUUUUU�?      �?                      �?;�;��?ى�؉��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?��K��K�?�����?�ǣ���?�+_�O�?�c�1��?�9�s��?�>�>��?[�[��?'u_[�?[4���?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?        d!Y�B�?�Mozӛ�?      �?        l�l��?��I��I�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�k(���?y�5���?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?                      �?�$I�$I�?n۶m۶�?d!Y�B�?�Mozӛ�?      �?      �?      �?                      �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?      �?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?              �?      �?        �������?�������?333333�?�������?      �?      �?              �?/�袋.�?F]t�E�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?�������?UUUUUU�?�q�q�?9��8���?�$I�$I�?n۶m۶�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        �{a���?GX�i���?7Āt,e�?��[��l�?�־a�?A��)A�?�x+�R�?:�&oe�?              �?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?        �-[�l��?ҤI�&M�?�袋.��?]t�E�?�?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��=���?a���{�?�.�袋�?F]t�E�?              �?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?	�=����?|a���?      �?        �������?�������?UUUUUU�?�������?              �?�q�q�?r�q��?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?              �?              �?        �t�bub��?     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ.s�ZhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�A         v       	          ����?�>�Ļ`�?9           ��@               /                    �?��,i��?           `{@                      
             �?Ɣ��Hr�?i             f@                                   �?Hm_!'1�?4            �X@                                 �_@t�6Z���?!            �K@       ������������������������       �                     ?@               
                    m@�q�q�?             8@              	       	          ����?؇���X�?
             ,@       ������������������������       �        	             (@        ������������������������       �                      @                                   �?���Q��?             $@                                  �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �E@               $                    �?�6i����?5            �S@                                  c@�?�P�a�?'             N@                                 `]@�Ń��̧?             E@                                   �?$�q-�?	             *@       ������������������������       �                     "@                                   \@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     =@                                  �g@�q�q�?             2@        ������������������������       �                     @                                   �?z�G�z�?
             .@                                  xq@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                !                   �^@ףp=
�?             $@        ������������������������       �                     @        "       #                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        %       &                    h@D�n�3�?             3@        ������������������������       �                     @        '       (                    �D@�n_Y�K�?
             *@        ������������������������       �                      @        )       .                    �?���!pc�?	             &@       *       -                    �?���Q��?             @       +       ,                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        0       k                    �?HO/�ն�?�            Pp@       1       H                    �?t�6Z���?�            �k@        2       ;       
             �?p���h�?@            @[@        3       :                   `n@�eP*L��?             &@       4       9                    @L@      �?              @       5       6                    �H@؇���X�?             @        ������������������������       �                     @        7       8                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        <       A                    �?`�(c�?9            �X@        =       >                    �?����X�?             @        ������������������������       �                     �?        ?       @                   �a@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        B       C                   Hp@@��,B�?4            �V@       ������������������������       �        !             L@        D       E       	          @33�?��?^�k�?            �A@       ������������������������       �                    �@@        F       G                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       d                   �c@���@��?J            �[@       J       S                     L@�E����?1             R@       K       P                   �b@�������?             F@       L       O       
             �?R���Q�?             D@        M       N       	          @33�?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �@@        Q       R                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        T       W                    �N@      �?             <@        U       V                   �e@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        X       c                    �?      �?             0@       Y       `                    �P@z�G�z�?             .@       Z       _                     P@�8��8��?             (@       [       \                    �O@r�q��?             @       ������������������������       �                     @        ]       ^                   @t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        a       b                   �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        e       j                    ]@ ���J��?            �C@        f       i                   �p@      �?              @        g       h                   p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ?@        l       s                    �?�p ��?            �D@        m       n                    �L@z�G�z�?
             .@       ������������������������       �                     $@        o       r                    �?���Q��?             @       p       q                    a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        t       u       
             �?�	j*D�?             :@       ������������������������       �        
             2@        ������������������������       �                      @        w       �                   �b@��*��?+            ~@       x       �                    �?�T|n�q�?�            0x@       y       �                   ``@�T`�[k�?�            �p@       z       �                    �?�gtq���?U            �`@        {       �                    �?      �?             L@        |       �       
             �?�q�q�?             ;@       }       �                    �O@8�A�0��?	             6@       ~       �       
             �?�E��ӭ�?             2@               �                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?������?             .@       �       �       	          033�?�	j*D�?             *@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       	             @J�8���?             =@       �       �                    �?�q�q�?             8@        ������������������������       �                     $@        �       �                   �]@X�Cc�?             ,@        ������������������������       �                      @        �       �                     M@      �?             (@       ������������������������       �                     @        �       �                   @_@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�6i����?8            �S@        �       �                    �H@X�<ݚ�?             "@        ������������������������       �                     @        �       �       	             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �Z@z��R[�?3            �Q@        �       �                   �o@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?���-T��?/             O@       �       �                    �L@h�WH��?'             K@       �       �                    \@$G$n��?            �B@        �       �                   �^@X�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @j@h�����?             <@       �       �                    @L@$�q-�?             *@       ������������������������       �        	             &@        �       �                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     1@        �       �                    �I@      �?              @        ������������������������       �                     �?        �       �                   `b@և���X�?             @       �       �       	          `ff�?���Q��?             @        ������������������������       �                      @        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �? ����?P            @`@       �       �       
             �?��4+̰�?;            @X@       �       �                    �?�E�����?5            �V@       ������������������������       �        '            �P@        �       �                   �e@�nkK�?             7@       ������������������������       �                     5@        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   Pv@����X�?             @       �       �       	             �?r�q��?             @       ������������������������       �                     @        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `a@�q�q�?            �@@        ������������������������       �                     &@        �       �       
             �?      �?             6@       �       �                   Pk@b�2�tk�?
             2@        �       �                     I@      �?              @        ������������������������       �                     �?        �       �                    �P@؇���X�?             @       �       �                   `c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �       
             �? ;=֦��?J            �^@        ������������������������       �                     ;@        �       �                   �Y@�==Q�P�?;            �W@        �       �                   @W@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                   pb@`��>�ϗ?3            @U@       ������������������������       �        %            �P@        �       �                    c@�}�+r��?             3@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        �             	          `ff@���3E��?<            @W@       �       �                    �?<�\`*��?7             U@        �       �                    �?l��
I��?             ;@        �       �       	          ����?��S���?	             .@       �       �                    \@z�G�z�?             $@        ������������������������       �                     @        �       �                    �F@�q�q�?             @        ������������������������       �                     �?        �       �                   pd@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@�8��8��?
             (@       �       �                    q@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�k�'7��?$            �L@        ������������������������       �                     5@        �       �                   �`@�E��ӭ�?             B@       �       �                   Pm@�C��2(�?             6@        �       �                   �\@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     &@        �                         f@և���X�?
             ,@       �                          �?�q�q�?             (@                                  b@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                    
             �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KMKK��hb�Bp  Qm4��?X��;�?�C2�<�?gx��m��?#h8����?��c+���?9/���?Y�Cc�?��)A��?X���oX�?              �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?        333333�?�������?�������?�������?      �?                      �?      �?                      �?kq�w��?T:�g *�?DDDDDD�?�����ݽ?��<��<�?�a�a�?�؉�؉�?;�;��?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?333333�?�������?      �?                      �?�������?�������?      �?        �������?�������?              �?      �?        (������?l(�����?              �?;�;��?ى�؉��?              �?F]t�E�?t�E]t�?�������?333333�?      �?      �?              �?      �?                      �?      �?        ��B�}��?�5��	��?X���oX�?��)A��?l�O����?�,�M�ɲ?t�E]t�?]t�E�?      �?      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?��)x9�?և���X�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?`��_���?h�h��?      �?        _�_��?�A�A�?      �?              �?      �?              �?      �?        L�Ϻ��?к����?r�q��?�q�q�?t�E]t�?/�袋.�?333333�?333333�?�$I�$I�?۶m۶m�?              �?      �?              �?              �?      �?              �?      �?              �?      �?UUUUUU�?�������?              �?      �?              �?      �?�������?�������?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?��-��-�?�A�A�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        8��18�?dp>�c�?�������?�������?      �?        �������?333333�?      �?      �?      �?                      �?      �?        ;�;��?vb'vb'�?              �?      �?        wwwwww�?""""""�?6eMYS��?���)k��?"5�x+��?���!5��?�\y@���?�Q�ߦ�?      �?      �?UUUUUU�?UUUUUU�?/�袋.�?颋.���?r�q��?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?�?wwwwww�?;�;��?vb'vb'�?      �?                      �?              �?      �?                      �?�rO#,��?|a���?UUUUUU�?�������?      �?        %I�$I��?�m۶m��?              �?      �?      �?      �?        �������?333333�?              �?      �?                      �?T:�g *�?kq�w��?r�q��?�q�q�?              �?�������?UUUUUU�?      �?                      �?X|�W|��?���?      �?      �?      �?                      �?�RJ)���?[k���Z�?B{	�%��?��^B{	�?���L�?к����?�q�q�?r�q��?              �?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?;�;��?�؉�؉�?              �?      �?      �?              �?      �?                      �?              �?      �?      �?      �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�����?�ȍ�ȍ�? tT����?_\����?l�l��?P��O���?              �?d!Y�B�?�Mozӛ�?              �?      �?      �?              �?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?9��8���?�8��8��?      �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?                      �?      �?        XG��).�?�%C��6�?              �?�a�+�?��%N��?�������?�������?              �?      �?        �?�������?              �?(�����?�5��P�?UUUUUU�?UUUUUU�?              �?      �?                      �?��.���?'�h��&�?=��<���?�a�a�?h/�����?Lh/����?�������?�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?-����b�?Lg1��t�?      �?        �q�q�?r�q��?]t�E�?F]t�E�?/�袋.�?F]t�E�?              �?      �?              �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?333333�?�������?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ8��`hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�E         �                    �?T �����??           ��@              [       
             �?��Z�b&�?L           ��@               $                    �?���g�?�            �i@                                  �L@>a�����?F            �Y@               
                    �? "��u�?#             I@                      	          ����?      �?             @        ������������������������       �                      @               	                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     F@                                  @R@      �?#             J@        ������������������������       �                     @                                   �?     ��?"             H@                                    N@���Q��?
             .@        ������������������������       �                     @                                  pc@      �?             (@                                 �`@"pc�
�?             &@                                  �?�q�q�?             @                                  �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?               #                   `@�C��2(�?            �@@              "                   �_@     ��?             0@                                   O@@4և���?             ,@       ������������������������       �                     "@               !                    �?z�G�z�?             @                                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        %       Z                    @R@�n_Y�K�?A             Z@       &       1       	          ����?���Q �??            �X@        '       .                     P@�q�q�?             8@       (       )       
             �?���N8�?             5@        ������������������������       �                      @        *       -                    �?�S����?             3@        +       ,                    �I@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             ,@        /       0                   Pa@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        2       M                    �?D˩�m��?.            �R@       3       H       	          `ff@�חF�P�?$             O@       4       ?                     N@4��?�?             J@       5       6                    �? �#�Ѵ�?            �E@        ������������������������       �        
             1@        7       8                    @I@$�q-�?             :@       ������������������������       �                     0@        9       :                    @J@z�G�z�?             $@        ������������������������       �                     �?        ;       <                   @q@�����H�?             "@        ������������������������       �                     @        =       >                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        @       A                    �?�q�q�?             "@        ������������������������       �                      @        B       C                   �`@؇���X�?             @        ������������������������       �                     @        D       G                    @      �?             @       E       F                    �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        I       L                   @n@      �?             $@       J       K                   0`@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        N       S                   �c@�q�q�?
             (@        O       P                   @l@r�q��?             @       ������������������������       �                     @        Q       R                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                    �H@�q�q�?             @        ������������������������       �                     �?        V       Y       	          033�?z�G�z�?             @        W       X                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        \       g                   @E@>4և�z�?�             u@        ]       f       	             �?�q�q�?             ;@       ^       c                   `@      �?             2@       _       `                   �_@���!pc�?             &@       ������������������������       �                     @        a       b                   �]@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        d       e                   @d@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        h       }                    �?���z�k�?�            Ps@        i       z       	          ����?
��[��?            @P@       j       y                   �c@d}h���?             L@       k       r                    �?H%u��?             I@        l       m                    �G@�n_Y�K�?             *@        ������������������������       �                     @        n       q                    �?�����H�?             "@        o       p                    �M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        s       x                    �?�?�|�?            �B@        t       u                    @L@��S�ۿ?             .@        ������������������������       �                     $@        v       w                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             6@        ������������������������       �                     @        {       |                    a@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ~       �                   @[@�2<�Z��?�            �n@               �                    �?�X����?             6@       �       �                    �J@�<ݚ�?	             2@       ������������������������       �                     (@        �       �                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �d@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   Pd@�v�ɱ?�            �k@       �       �                    @�}�+r��?]             c@       �       �       	          ����?˒�#�?Y            �b@       �       �                    @L@@ݚ)�?V             b@       ������������������������       �        G            �]@        �       �                   @t@���B���?             :@       �       �                    �?�J�4�?             9@       �       �                    b@z�G�z�?
             4@       �       �                   Hp@�����H�?	             2@       ������������������������       �                     (@        �       �       	          @33�?�q�q�?             @        ������������������������       �                     @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   h@      �?             @        ������������������������       �                      @        �       �                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        +            �Q@        �       �       
             �?PcG���?�            �w@       �       �                    �?�ţ����?�            0t@        �       �       
             �?r٣����?            �@@        �       �                    �I@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@�+$�jP�?             ;@       �       �                    �?     ��?             0@       �       �                   xt@�n_Y�K�?             *@       �       �                   �a@���!pc�?
             &@       �       �                    �M@      �?              @       ������������������������       �                     @        �       �                     O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Hp@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             &@        �       �                   �[@�������?�             r@        �       �                    �?f���M�?             ?@        �       �       	          ����?      �?              @        �       �       	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?��<b���?             7@        ������������������������       �                     "@        �       �                     N@X�Cc�?	             ,@       �       �                   @Y@      �?             $@        ������������������������       �                     @        �       �       
             �?����X�?             @        ������������������������       �                     @        �       �                    �K@      �?             @       �       �                   �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �R@���VҴ?�            0p@       �       �                   �e@ �?�            �o@       �       �                   �b@������?�            �o@       �       �       	          ���@Pl0�ͤ?�             n@       �       �                    @L@ �LV�-�?�            �j@        ������������������������       �        ?             Y@        �       �                    �?��x$�?G            �\@       �       �                   `Z@��<b�ƥ?9             W@        �       �                   0g@$�q-�?             :@        ������������������������       �                     *@        �       �                   �W@8�Z$���?	             *@        ������������������������       �                     @        �       �                   Pk@����X�?             @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   `a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        (            �P@        �       �                    �?�nkK�?             7@       ������������������������       �                     3@        �       �                   0`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   p@$�q-�?             :@       ������������������������       �                     4@        �       �                    `@�q�q�?             @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	             �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                   @`@�q�q�?             @        ������������������������       �                     �?        �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                         Pj@~|z����?$            �J@        �                         @b@�q�q�?             8@       �                         @e@r�q��?             2@       �                          �?�t����?             1@       �                         `b@"pc�
�?             &@       �                           P@���Q��?             @       �                           I@�q�q�?             @       �       �                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?                                 �N@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        	                          K@����"�?             =@        
                         o@r�q��?
             (@       ������������������������       �                     "@                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                hp@��.k���?             1@                                @a@z�G�z�?             $@                               �`@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                xt@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�Bp  ��G��G�?�\�\�?�h_����?J.A�~��?C����?^�	���?�?�������?���Q��?�G�z�?      �?      �?              �?      �?      �?      �?                      �?              �?      �?      �?      �?              �?      �?�������?333333�?      �?              �?      �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        F]t�E�?]t�E�?      �?      �?�$I�$I�?n۶m۶�?              �?�������?�������?      �?      �?      �?                      �?              �?      �?                      �?;�;��?ى�؉��?9/����?����>4�?�������?�������?��y��y�?�a�a�?      �?        ^Cy�5�?(������?333333�?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        a�|���?}���g�?�Zk����?��RJ)��?�N��N��?ى�؉��?�/����?�}A_Ч?      �?        �؉�؉�?;�;��?      �?        �������?�������?              �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?      �?              �?      �?              �?              �?      �?UUUUUU�?�������?      �?                      �?      �?        �������?�������?UUUUUU�?�������?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?      �?              �?      �?              �?                      �?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?t�E]t�?F]t�E�?              �?333333�?�������?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?              �?���O ��?ch���V�?7r#7r#�?�����?I�$I�$�?۶m۶m�?)\���(�?���Q��?;�;��?ى�؉��?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        *�Y7�"�?к����?�������?�?      �?        �������?�������?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?              �?      �?        mާ�d�?.�u�y�?�E]t��?]t�E]�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?        ��w����?5'��Ps�?�5��P�?(�����?�g�`�|�?v�)�Y7�?9��8���?r�qǡ?      �?        ��؉���?ى�؉��?�z�G��?{�G�z�?�������?�������?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?      �?              �?      �?              �?      �?      �?              �?      �?      �?                      �?      �?        br1��?}g���Q�?3@%[�Ʒ?�W�"�?|���?>���>�?      �?      �?      �?                      �?B{	�%��?/�����?      �?      �?ى�؉��?;�;��?t�E]t�?F]t�E�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?%�6Q�k�?�(ٵ���?��Zk���?��RJ)��?      �?      �?      �?      �?      �?                      �?      �?        ��Moz��?��,d!�?              �?�m۶m��?%I�$I��?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�[�þ�?A����?�?�������?�q�q�?�q�q�?�>�>�?�
V�
V�?X:Ɂ���?��i���?              �?��s���?�aܯK*�?d!Y�B�?��7��M�?;�;��?�؉�؉�?              �?;�;��?;�;��?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?d!Y�B�?�Mozӛ�?              �?      �?      �?              �?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?/�袋.�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?        ��sHM0�?�	�[���?�������?�������?UUUUUU�?�������?�?<<<<<<�?F]t�E�?/�袋.�?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?              �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?	�=����?�i��F�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�?�������?�������?�������?�������?333333�?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�>�&hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK�h��B@<         d                   �`@�ʻ����?F           ��@               U                    �?��`�+"�?           z@              (                    �?�����?�            @r@                                   U@�ǧ\�?I            �Z@        ������������������������       �                     @                                   �?��ȯ��?F            �Y@                      	          433�?      �?             @@              	                    �?���7�?             6@       ������������������������       �                     4@        
                           @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?�z�G��?             $@                                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?              @                                 �n@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?               #                    �?��(@��?/            �Q@                     
             �?T�7�s��?&            �L@                      	             �?(;L]n�?             >@                                 �Y@�IєX�?
             1@        ������������������������       �                     �?        ������������������������       �        	             0@        ������������������������       �        	             *@               "                   @c@�����H�?             ;@                                   �?�q�q�?             "@        ������������������������       �                     �?                !                   @_@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        $       '                   �^@$�q-�?	             *@        %       &       	          @33�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        )       4                    �?d�J U��?y            @g@        *       +                   �Z@X�Cc�?
             ,@        ������������������������       �                     @        ,       1                    �?����X�?             @       -       .                   �`@z�G�z�?             @        ������������������������       �                      @        /       0       	            �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        2       3                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       T                    �M@ �#�Ѵ�?o            �e@       6       9                    [@���l��?G            �[@        7       8                    �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        :       S                    @HQ˄�ľ?E            @[@       ;       L                    �?�X�<ݺ?D             [@       <       A                    @L@X;��?8            @V@       =       @       	             �?�k~X��?-             R@        >       ?                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        &             P@        B       C                    �?�t����?             1@        ������������������������       �                     @        D       K                   �r@z�G�z�?             $@       E       F       
             �?�����H�?             "@        ������������������������       �                      @        G       J                     M@؇���X�?             @       H       I                   @[@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        M       R       	             @�S����?             3@       N       Q                   �Z@�IєX�?             1@        O       P                    @K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        (            �N@        V       ]                     Q@0{�v��?M            @_@       W       X       
             �?����q�?D            @[@       ������������������������       �        9            @V@        Y       Z                    \@ףp=
�?             4@       ������������������������       �                     .@        [       \                     O@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ^       _                    �?     ��?	             0@        ������������������������       �                      @        `       a                   c@X�Cc�?             ,@       ������������������������       �                     @        b       c                   �[@      �?              @        ������������������������       �                     @        ������������������������       �                     @        e       �                    �?��Q/��?7           P@       f       �                    �?p6��%�?�            �x@       g       �       
             �?��%c�?�            �t@        h       �                   `a@��9܂�?4            @V@       i       �       	             @������?'            @Q@       j       }                   q@     8�?#             P@       k       l                    T@�J��%�?            �H@        ������������������������       �                     @        m       n                    �?      �?             F@        ������������������������       �        	             4@        o       p                   �a@r�q��?             8@        ������������������������       �                     @        q       |                    �L@�����?             3@       r       {                    @L@      �?	             (@       s       t                    �?���Q��?             $@        ������������������������       �                      @        u       v                    �?      �?              @        ������������������������       �                      @        w       x                   @b@�q�q�?             @        ������������������������       �                      @        y       z                    �J@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ~       �                   �e@������?             .@              �                     O@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �l@ףp=
�?             4@        �       �                    @      �?             @        ������������������������       �                      @        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �e@      �?	             0@       ������������������������       �                     .@        ������������������������       �                     �?        �       �       	          033@�1~�?�            `n@       �       �                    �L@���i��?�             n@       �       �                   0h@ f^8���?}            �i@       �       �                   `\@p7 .���?{            `i@        �       �                    �?�J�4�?             9@       �       �                   d@"pc�
�?             6@       �       �                   �b@�	j*D�?	             *@       ������������������������       �                      @        �       �                    �J@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                   �f@@~��?i            @f@       ������������������������       �        ]             d@        �       �                   �f@�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �                     1@        �       �                   �h@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0c@4�2%ޑ�?            �A@       �       �                    ]@      �?             0@        �       �                   @n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                   �`@p�ݯ��?             3@        ������������������������       �                     @        �       �                    s@؇���X�?             ,@       �       �                    b@$�q-�?             *@       ������������������������       �                     "@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?N1���?(            �N@        �       �       
             �?��s����?             5@        ������������������������       �                     "@        �       �                   @[@�q�q�?	             (@       ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?���Q��?             D@        �       �       
             �?ҳ�wY;�?             1@        ������������������������       �                      @        �       �                   ``@������?
             .@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   @c@�q�q�?             @        ������������������������       �                     �?        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@ףp=
�?             $@       �       �                   q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   0a@��<b���?             7@        �       �                   �`@X�Cc�?             ,@       �       �                    �L@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�<ݚ�?F             [@       �       �                   Pd@�:�^���?3            �S@       �       �                   �Z@Х-��ٹ?1            �R@        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    a@������?/             R@       ������������������������       �                    �B@        �       �                    �M@ >�֕�?            �A@       �       �                   `a@ףp=
�?             4@        ������������������������       �                     �?        �       �                     M@�}�+r��?             3@       ������������������������       �        
             .@        �       �                   �b@      �?             @        ������������������������       �                      @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             .@        ������������������������       �                     @        �       �                    f@*;L]n�?             >@       �       �                   �b@$��m��?             :@       �       �                    �?X�Cc�?
             ,@        ������������������������       �                     �?        �       �                    �?�	j*D�?	             *@       �       �                   pa@���Q��?             $@        ������������������������       �                      @        �       �                   �[@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  <<<<<<�?�������?��<}��?�Eΰ�R�?�#F��?<w�ܹs�?�&oe��?���!5��?              �?dddddd�?777777�?      �?      �?�.�袋�?F]t�E�?      �?              �?      �?      �?                      �?ffffff�?333333�?      �?      �?              �?      �?              �?      �?�m۶m��?�$I�$I�?      �?                      �?      �?        ����?��+��+�?�}��?p�}��?�?�������?�?�?      �?                      �?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        �؉�؉�?;�;��?�������?�������?      �?                      �?      �?        �Gy�?�7�p��?�m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�}A_Ч?�/����?5'��Ps�?��蕱�?      �?      �?              �?      �?        ��p�?߅����?�q�q�?��8��8�?�E(B�?�u�{���?�q�q�?�8��8��?      �?      �?      �?                      �?              �?�?<<<<<<�?              �?�������?�������?�q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?        ^Cy�5�?(������?�?�?      �?      �?              �?      �?                      �?      �?              �?                      �?;�O��n�?V-��?�,�M�ɒ?���%�i�?              �?�������?�������?              �?�������?333333�?      �?                      �?      �?      �?      �?        �m۶m��?%I�$I��?              �?      �?      �?              �?      �?        �-Nk�O�?�c)�`�?��0�]��?BJ�eD�?.+Jx��?GS��r�?�.p��? ��G?��??���(�?ہ�v`��?     ��?      �?c}h���?9/����?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?Q^Cy��?^Cy�5�?      �?      �?333333�?�������?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �?wwwwww�?;�;��?;�;��?              �?      �?              �?                      �?�������?�������?      �?      �?              �?      �?      �?              �?      �?              �?      �?              �?      �?        -����?�F�� ۰?�$�$�?$�$��?H%�e�?��VCӝ?Ŭ�:6�?igJ��8�?�z�G��?{�G�z�?/�袋.�?F]t�E�?vb'vb'�?;�;��?      �?        �������?�������?              �?      �?              �?              �?        ��G?���?p�\�w?      �?        ��8��8�?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�A�A�?      �?      �?      �?      �?      �?                      �?      �?        ^Cy�5�?Cy�5��?              �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?      �?              �?      �?              �?      �?                      �?              �?�}�K�`�?�:ڼO�?�a�a�?z��y���?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?�������?�������?      �?        �?wwwwww�?333333�?�������?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?��,d!�?��Moz��?%I�$I��?�m۶m��?/�袋.�?F]t�E�?      �?                      �?              �?      �?        �q�q�?9��8���?�o��o��?� � �?O贁N�?K~��K�?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?�A�A�?��+��+�?�������?�������?      �?        (�����?�5��P�?              �?      �?      �?              �?      �?      �?      �?                      �?              �?      �?        """"""�?�������?�N��N��?vb'vb'�?�m۶m��?%I�$I��?      �?        ;�;��?vb'vb'�?�������?333333�?      �?              �?      �?      �?                      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�w}@hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@F         �                    �?�LT ���?D           ��@                                 �_@��CU�G�?;           0@                                  �U@�.ߴ#�?O            �^@        ������������������������       �                     �?                      
             �?���tcH�?N            @^@       ������������������������       �        :             W@                                   �?д>��C�?             =@        ������������������������       �                     �?        	       
                    �?�>4և��?             <@        ������������������������       �                     �?                                   @M@�+$�jP�?             ;@                                  �?�IєX�?             1@                     	          ����?�C��2(�?             &@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  �b@���Q��?             $@                                 �_@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @               �                    �?������?�            �w@              n       
             �?�Xp��?�             s@              G       	             �?#n��?            �j@               @                   �b@�	j*D�?3            �V@              !                    �?DE��2{�?+            �R@                                    �?�����H�?             "@                                  �p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        "       #       	          ����?�GN�z�?$            �P@        ������������������������       �                     3@        $       ?                   �a@(���@��?            �G@       %       8                    �?�Gi����?            �B@       &       '                   �g@���@M^�?             ?@        ������������������������       �                      @        (       3                    @M@
;&����?             7@       )       *                   �l@j���� �?	             1@        ������������������������       �                     @        +       2                    a@�q�q�?             (@       ,       -       	          433�?      �?              @        ������������������������       �                     �?        .       1                    @J@����X�?             @       /       0                   �t@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        4       5                   �o@�q�q�?             @        ������������������������       �                      @        6       7                   p`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        9       :                    �I@      �?             @        ������������������������       �                      @        ;       <                   `Z@      �?             @        ������������������������       �                      @        =       >                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        A       F       	          @33�?      �?             0@       B       E                    �J@X�<ݚ�?             "@       C       D                   ``@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        H       I                   �Z@�7���?L             _@        ������������������������       �                      @        J       W                    �?�٠n�}�?K            �^@        K       L                   �c@      �?             0@        ������������������������       �                      @        M       N       
             �?؇���X�?
             ,@        ������������������������       �                      @        O       R                    �?r�q��?	             (@        P       Q                    �O@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        S       V                    �J@؇���X�?             @        T       U                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        X       c       	          ����?����?@            �Z@        Y       Z       
             �?ܷ��?��?             =@        ������������������������       �                     @        [       b                    �?�LQ�1	�?             7@       \       ]                    �G@r�q��?	             2@        ������������������������       �                      @        ^       a                   �i@      �?             0@        _       `                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     @        d       i                    _@�g<a�?2            @S@        e       f       	          033@@4և���?
             ,@       ������������������������       �                     (@        g       h                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        j       k                   q@ ������?(            �O@       ������������������������       �                     G@        l       m                   �q@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@        o       �                    @O@:��?:            @V@       p                           �?�(�Tw��?2            �S@        q       z                   �_@�eP*L��?             6@       r       s                    �?      �?             (@        ������������������������       �                     �?        t       u                   �^@"pc�
�?             &@        ������������������������       �                     �?        v       w                    �G@ףp=
�?             $@       ������������������������       �                     @        x       y                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        {       ~       	             �?�z�G��?             $@       |       }                     N@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �I@�>4և��?#             L@       �       �       	          433�?@4և���?             <@       �       �                   pf@`2U0*��?             9@       ������������������������       �                     8@        ������������������������       �                     �?        �       �                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @J@����X�?             <@        ������������������������       �                      @        �       �                    @K@�θ�?             :@        ������������������������       �                     @        �       �                    @N@����X�?             5@       �       �       	          033�?�q�q�?	             .@       �       �       	          ����?r�q��?             (@       �       �                    �?ףp=
�?             $@       �       �                   �b@�q�q�?             @        ������������������������       �                     �?        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                   �k@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@���!pc�?             &@       �       �                    [@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?L������?3            @R@       �       �                    �R@      �?,             P@       ������������������������       �        +             O@        ������������������������       �                      @        �       �                   �l@�q�q�?             "@        ������������������������       �                     @        �       �                    �G@      �?             @        ������������������������       �                      @        �       �                    Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?�	�lW��?	           0z@       �       �       
             �?fe�07�?�            �q@        �       �                    �?����5�?$            �N@       �       �                    �?\X��t�?             G@        �       �                   �q@ҳ�wY;�?
             1@       �       �                    �?�8��8��?             (@        �       �                    �J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?8^s]e�?             =@       �       �                    �J@8�A�0��?             6@        ������������������������       �                      @        �       �       	          ����?X�Cc�?             ,@       �       �                    �L@X�<ݚ�?             "@       �       �                   �p@�q�q�?             @       �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             .@        �       �                   @n@ �Jj�G�?�            �k@       ������������������������       �        T            ``@        �       �                   0c@ p�/��?<            @V@        �       �                    �M@������?            �B@       �       �                   �b@؇���X�?             <@       �       �                    �?$�q-�?             :@        �       �                     @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     L@�nkK�?             7@       ������������������������       �                     2@        �       �                   �_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �        "             J@        �             
             �?ڡ�:x��?U            @a@       �       �                    �B@     ��?=             X@        �       �                   (p@����X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �                          �?�)V���?9            @V@        �       �                    @�>$�*��?            �D@       �       �                    �?���|���?            �@@        �       �                    c@      �?              @       �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?`�Q��?             9@       �       �                   �c@���N8�?             5@       �       �       	          `ff�?r�q��?
             2@        �       �                    �?և���X�?             @       �       �                   `Z@�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       	             @      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �                           X@      �?              @        ������������������������       �                     �?                                  P@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                �\@8��8���?             H@        ������������������������       �                     @                                �`@t��ճC�?             F@       ������������������������       �                     <@                                 �?     ��?	             0@       	      
                   �?@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                      @                                �]@r�q��?             E@                                Pa@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �L@�?�'�@�?             C@       ������������������������       �                     6@                                 @O@     ��?
             0@                               �a@      �?              @        ������������������������       �                     @        ������������������������       �                     @                                 �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �t�b��7     h�h)h,K ��h.��R�(KMKK��hb�B�  ��u���?�(E~��?8��ѽ��?���P��?XG��).�?�K�`m�?      �?        �C��2(�?����|��?              �?|a���?a���{�?              �?�m۶m��?�$I�$I�?              �?B{	�%��?/�����?�?�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�������?333333�?�$I�$I�?۶m۶m�?      �?                      �?      �?        ��3T���?@2�խ �?�k(���?��k(��?hsy�7�?& �a2�?;�;��?vb'vb'�?O贁N�?,�Œ_,�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E�?�袋.��?              �?R�٨�l�?W�+���?#�u�)��?o0E>��?�c�1��?�s�9��?              �?Y�B��?�Mozӛ�?�������?ZZZZZZ�?      �?        �������?�������?      �?      �?              �?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?              �?      �?      �?r�q��?�q�q�?۶m۶m�?�$I�$I�?              �?      �?              �?              �?        ��Zk���?)��RJ)�?      �?        �u�y��?Pq����?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?�������?�������?�������?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?�V�9�&�?��`��}�?a���{�?��=���?              �?Y�B��?��Moz��?UUUUUU�?�������?      �?              �?      �?      �?      �?              �?      �?                      �?              �?�cj`?���8+�?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?        AA�?��}��}�?              �?�?�?      �?                      �?S��Ԧ6�?Y�JV���?�o��o��?� � �?]t�E�?t�E]t�?      �?      �?      �?        F]t�E�?/�袋.�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?ffffff�?333333�?      �?      �?      �?                      �?              �?�$I�$I�?�m۶m��?n۶m۶�?�$I�$I�?���Q��?{�G�z�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?              �?ى�؉��?�؉�؉�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?�������?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?              �?      �?              �?      �?                      �?�������?UUUUUU�?      �?              �?      �?              �?      �?        t�E]t�?F]t�E�?�q�q�?�q�q�?      �?                      �?      �?        ����?�Ǐ?~�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?      �?                      �?������?���?��,'��?pMc��?������?��).��?��Moz��?!Y�B�?�������?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?	�=����?|a���?/�袋.�?颋.���?              �?%I�$I��?�m۶m��?�q�q�?r�q��?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?              �?      �?                      �?              �?k߰�k�?��)A��?      �?        �G?�я�?p�\��?��g�`��?к����?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�Mozӛ�?d!Y�B�?      �?        �������?�������?              �?      �?                      �?      �?              �?        �g��%�?̵s��?      �?      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?         ��G?��?p�\��?�����?�18���?F]t�E�?]t�E]�?      �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?{�G�z�?��(\���?��y��y�?�a�a�?UUUUUU�?�������?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?                      �?�������?UUUUUU�?      �?        t�E]t�?�E]t��?              �?      �?      �?�$I�$I�?n۶m۶�?      �?                      �?      �?        �������?UUUUUU�?      �?      �?              �?      �?        ������?y�5���?      �?              �?      �?      �?      �?              �?      �?              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJudxhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK酔h��B@:         n       	          ����?z�ГPo�?>           ��@               5                    �?�)s�Z�?           �|@                      
             �?�-ῃ�?n            �f@                                 �b@,�T�6�?<             Z@                     	          833�? �\���?/            �S@       ������������������������       �        (            �Q@                                   �?X�<ݚ�?             "@        ������������������������       �                     @        	       
                   �`@r�q��?             @       ������������������������       �                     @                                   b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �L@ �o_��?             9@                     	          833�?؇���X�?             5@                                  �?�IєX�?	             1@       ������������������������       �                     0@        ������������������������       �                     �?                                  ``@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  @E@�2��?2            �S@                                   a@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @                                    B@&�a2o��?,            @Q@        ������������������������       �                     @               "                    c@     8�?+             P@              !                    �?������?             B@                                    �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �@@        #       2                    �L@X�Cc�?             <@       $       +                   `\@�GN�z�?             6@        %       &                    �?և���X�?             @        ������������������������       �                     �?        '       (                    �?�q�q�?             @        ������������������������       �                     @        )       *                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ,       1                    �?��S�ۿ?	             .@       -       .                    �?ףp=
�?             $@        ������������������������       �                     @        /       0                   pf@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        3       4                   �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        6       Q       
             �?��K�"�?�            �q@        7       >                    �?�q�q�?,             R@        8       9                     G@������?             .@        ������������������������       �                     "@        :       =       	          ����?�q�q�?             @       ;       <                     P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ?       L                   0a@�k�'7��?             �L@       @       G       	          ����?��H�}�?             9@       A       F                    @J@      �?             0@        B       E                    f@�q�q�?             @       C       D                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        H       K                   Pm@�<ݚ�?             "@        I       J                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        M       N                     Q@      �?             @@       ������������������������       �                     >@        O       P                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        R       g                    �O@������?�             j@       S       `                    c@`��Zש?}             h@       T       ]       	            �?�h%�M��?p            `e@       U       V                    �?�������?l            �d@       ������������������������       �        E             \@        W       \                    �G@@3����?'             K@        X       [                   @[@ ��WV�?             :@        Y       Z                    @E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     <@        ^       _                     L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        a       f                   �d@��2(&�?             6@       b       e                   p@���!pc�?             &@       c       d                   pd@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        h       m       	          ����?���Q��?             .@       i       j                    `P@�eP*L��?             &@        ������������������������       �                     @        k       l                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        o       �                    _@�����?           p|@        p       �                    �?�ꮃG�?T            @a@       q       r                   ``@և���X�?+            �Q@        ������������������������       �                     .@        s       t                    �?���!pc�?            �K@        ������������������������       �                     .@        u       v                    `@      �?             D@        ������������������������       �                      @        w       |                    �?     ��?             @@        x       {                   Pd@      �?             @       y       z                    a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        }       �                   �d@8�Z$���?             :@       ~       �                    @�KM�]�?	             3@              �                    @B@r�q��?             (@        ������������������������       �                     �?        �       �                   �i@�C��2(�?             &@        �       �                   @g@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   m@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          033@�����?)             Q@       �       �                    �?(2��R�?#            �M@       �       �       
             �?p���?             I@        �       �                   �W@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     C@        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                   �\@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   pk@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?H��w&��?�            �s@       �       �                    @B@�1�`jg�?�            �k@        ������������������������       �                      @        �       �                    c@ '��h�?�            @k@       �       �       
             �?����?�            @i@       �       �                    �D@ ������?u            �g@        �       �       	             �?r�q��?             @       �       �                    _@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �? h'M#�?r            �f@        �       �                   `U@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        �       �                    @L@�=
ףp�?d             d@        ������������������������       �        1            @T@        �       �                   �`@�Fǌ��?3            �S@        �       �                    �L@$�q-�?	             *@        �       �                    e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �        *            �P@        �       �                   �`@8�Z$���?             *@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?     ��?
             0@       �       �                   �`@X�Cc�?             ,@        ������������������������       �                      @        �       �                    �?�q�q�?             (@        �       �                    �?r�q��?             @       �       �       	          ���@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                     P@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�U�!��?@            @X@        �       �                    \@�C��2(�?             6@        ������������������������       �                      @        ������������������������       �                     4@        �       �       	          pff�?X���[�?1            �R@        �       �                    �N@p�ݯ��?             C@       �       �       
             �?V�a�� �?             =@        �       �                    b@X�Cc�?	             ,@       �       �       	             �?X�<ݚ�?             "@       �       �                     I@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @��S�ۿ?	             .@       ������������������������       �                     &@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�����H�?             "@       �       �                   �c@r�q��?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �c@$G$n��?            �B@       �       �       
             �? 7���B�?             ;@        �       �       	          033@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     8@        �       �                   0e@���Q��?             $@        ������������������������       �                     @        �       �                   ``@؇���X�?             @       �       �                   �f@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  1�i�M��?��<Y �?SGQ��?Yq]�3��?�����?�).�u�?;�;��?ى�؉��?�3���?���7a�?              �?�q�q�?r�q��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�Q����?
ףp=
�?�$I�$I�?۶m۶m�?�?�?              �?      �?              �?      �?              �?      �?              �?        ���JG�?�&��jq�?�������?�������?              �?      �?        ��Q�g��?ہ�v`��?              �?     ��?      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        %I�$I��?�m۶m��?�袋.��?]t�E�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�?�������?�������?      �?        �������?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?              �?      �?        ����?|�W|�W�?�������?�������?wwwwww�?�?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?        Lg1��t�?-����b�?
ףp=
�?{�G�z�?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?                      �?9��8���?�q�q�?333333�?�������?      �?                      �?      �?              �?      �?              �?      �?      �?              �?      �?        ��N��N�?;�;��?aw&��+�?�1�K��?��/��?@��?(፦��?��k��x?      �?        ���Kh�?h/�����?O��N���?;�;��?      �?      �?      �?                      �?      �?              �?        �������?�������?      �?                      �?��.���?t�E]t�?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?                      �?              �?      �?        333333�?�������?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?                      �?      �?        � 	� 	�?�����?��Q�g��?;0�̵�?�$I�$I�?۶m۶m�?              �?F]t�E�?t�E]t�?      �?              �?      �?              �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?        ;�;��?;�;��?�k(���?(�����?�������?UUUUUU�?              �?]t�E�?F]t�E�?�������?�������?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?              �?      �?        xxxxxx�?�������?'u_[�?=�"h8��?{�G�z�?\���(\�?UUUUUU�?UUUUUU�?      �?                      �?              �?9��8���?�q�q�?      �?                      �?r�q��?�q�q�?      �?        �������?�������?      �?                      �?K_R����?-hk���?�־a�?A��)A�?      �?        �w� z|�?���]8��?z��~�X�?|#
L:5�?AA�?��}��}�?UUUUUU�?�������?      �?      �?              �?      �?                      �?�"Qj�a�?t�VNx��?d!Y�B�?�Mozӛ�?      �?                      �?������y?�������?              �?�3���?1���M��?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?              �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�m۶m��?%I�$I��?              �?�������?�������?UUUUUU�?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?���:*�? tT����?]t�E�?F]t�E�?              �?      �?        �X�%��?��:m��?^Cy�5�?Cy�5��?��{a�?a���{�?%I�$I��?�m۶m��?�q�q�?r�q��?�������?�������?              �?      �?                      �?      �?        �������?�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?���L�?к����?h/�����?	�%����?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?333333�?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJD ?<hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKم�h��B@6         n                    �?n�A��?=           ��@              1       
             �?Ds\�A�?W           Ѐ@                                   �?P�|

��?�             h@                                   b@��V#�?            �E@                     
             �?tk~X��?             B@        ������������������������       �                     @                                  �Q@<���D�?            �@@        ������������������������       �                      @        	       
                    �?`Jj��?             ?@       ������������������������       �                     =@        ������������������������       �                      @        ������������������������       �                     @               0                   �f@r�q��?f            �b@              !                   �l@x�5?,R�?b             b@                     	          ����?DE�SA_�?@            @X@        ������������������������       �                     E@                                    �O@t�6Z���?#            �K@                                  @O@� ��1�?            �D@                     
             �?������?            �B@                      	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                  �c@�FVQ&�?            �@@                                  @G@�g�y��?             ?@                                  �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     <@                                   �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             ,@        "       %       
             �?��|�5��?"            �G@        #       $       	          033@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        &       '                    _@      �?             D@        ������������������������       �        
             .@        (       /                   0o@z�G�z�?             9@        )       *                    �?      �?              @        ������������������������       �                     @        +       .                     N@���Q��?             @       ,       -                    @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     @        2       m       	          ���@0��a�?�            �u@       3       @                    P@�Yr8{�?�            pu@        4       5                   `X@���>4��?             <@        ������������������������       �                     @        6       7                   �^@\X��t�?             7@        ������������������������       �                     @        8       =                    �?j���� �?             1@       9       <                   �b@      �?              @       :       ;                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        >       ?                   �a@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        A       l                   @g@��S�ۿ?�            �s@       B       Y                    �?�U��w1�?�            �s@        C       H                   �a@�M���?.             Q@       D       E       	             �?      �?             @@       ������������������������       �                     >@        F       G                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       N                   @^@b�2�tk�?             B@        J       M                   Pl@�q�q�?             .@        K       L                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        O       T                    b@��s����?             5@       P       Q                     L@      �?             0@       ������������������������       �                      @        R       S                   �q@      �?              @        ������������������������       �                     @        ������������������������       �                      @        U       X                   �d@���Q��?             @       V       W                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        Z       e                    @ �ƭr�?�            �n@       [       \                    @L@�H�I���?�            @l@       ������������������������       �        p            �g@        ]       b                   ht@@-�_ .�?            �B@       ^       a                    �L@Pa�	�?            �@@        _       `                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     >@        c       d                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        f       k                   a@�KM�]�?             3@        g       h                    h@�q�q�?             @        ������������������������       �                      @        i       j                   �j@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                      @        o       �       
             �?�"�q��?�            �w@       p       s                   �Z@���R���?�            �s@        q       r                   0a@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        t       �                    �?��7H�?�            ps@       u       �                    �?������?�            `n@       v       �                   �b@����\�?j            �f@       w       �       	          ����?x%�%%ն?e            `e@       x       �                    �L@��y� �?6            @W@       y       �                    @K@L紂P�?!            �I@       z       {                   pb@�}�+r��?             C@       ������������������������       �                     :@        |                          `c@r�q��?             (@        }       ~                   @\@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �K@�n_Y�K�?	             *@        �       �                   0p@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�z�G��?             $@       ������������������������       �                     @        �       �                   @_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �O@�Ń��̧?             E@       ������������������������       �                     :@        �       �                    �?      �?             0@       �       �                   �`@�C��2(�?             &@        �       �                   p`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �        /            �S@        �       �       	          433�?�q�q�?             "@        ������������������������       �                     @        �       �                   �c@      �?             @       �       �                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @s@���N8�?+            �O@       ������������������������       �        %            �J@        �       �                    �?�z�G��?             $@        ������������������������       �                     @        �       �       
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@������?'             Q@       �       �                    �?�Ń��̧?             E@        �       �                   �Z@�����H�?             "@       ������������������������       �                     @        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �@@        �       �                    �?
j*D>�?             :@       �       �       	             �?      �?             6@        ������������������������       �                     @        �       �                    �?D�n�3�?             3@        ������������������������       �                     @        �       �                   �\@��S���?	             .@        ������������������������       �                     �?        �       �                   �l@և���X�?             ,@        �       �       	             �?r�q��?             @       �       �                   c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    n@      �?              @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�g�y��?%             O@       �       �                   `b@v�X��?             F@       �       �       	          ����?���@��?            �B@        �       �                    �?�q�q�?             "@       �       �                   @`@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@4և���?             <@       �       �       	          033�?�����?             5@       ������������������������       �                     2@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �M@����X�?             @       �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�X�<ݺ?
             2@       ������������������������       �                     .@        �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  >��=���?a�a��?�0���x�?�}lF�?n����?I	9��?eMYS֔�?6eMYS��?r�q��?9��8���?              �?|���?|���?              �?���{��?�B!��?      �?                      �?              �?UUUUUU�?�������?9��8���?r�q��?����?���_\�?              �?��)A��?X���oX�?������?������?к����?��g�`��?      �?      �?      �?                      �?|���?>����?�B!��?��{���?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?      �?                      �?x6�;��?br1���?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?              �?�������?�������?      �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �+MX�y�?á�=u2�?�L��2��?���i޺?n۶m۶�?I�$I�$�?              �?!Y�B�?��Moz��?      �?        ZZZZZZ�?�������?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?      �?        r�q��?�q�q�?      �?                      �?�������?�?�^�׸�?�:�r�?�������?<<<<<<�?      �?      �?      �?              �?      �?              �?      �?        �8��8��?9��8���?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?z��y���?�a�a�?      �?      �?      �?              �?      �?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        Ӟ�@z�?ȝ%�淐?x�!���?x�!���?      �?        S�n0E�?к����?|���?|���?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�k(���?(�����?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?                      �?              �?|n�S���?a�+F�?2��X��?J�-�?�m۶m��?�$I�$I�?              �?      �?        �Σ�)�?,�����?�:���?�������?�>�>�?.؂-؂�?@���?�/����?X`��??���O?�?�������?�������?(�����?�5��P�?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?ى�؉��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?333333�?ffffff�?              �?      �?      �?              �?      �?        �a�a�?��<��<�?              �?      �?      �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?      �?              �?      �?                      �?�a�a�?��y��y�?              �?333333�?ffffff�?              �?      �?      �?      �?                      �?�?xxxxxx�?�a�a�?��<��<�?�q�q�?�q�q�?              �?      �?      �?              �?      �?                      �?b'vb'v�?;�;��?      �?      �?              �?l(�����?(������?      �?        �������?�?      �?        ۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        ��{���?�B!��?颋.���?�.�袋�?к����?L�Ϻ��?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?              �?      �?              �?      �?              �?      �?        �$I�$I�?n۶m۶�?�a�a�?=��<���?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��UhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�=         �       
             �?�HK��x�??           ��@              W                    �?� �(���?Q           Ѐ@                                  �? w�����?�            pw@                                  pm@�����?            �H@        ������������������������       �        
             4@                                  pn@J�8���?             =@        ������������������������       �                     @                                  �r@R�}e�.�?             :@        	       
                    �H@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@                                   b@���Q��?             .@                                  y@�q�q�?             @                                 �`@z�G�z�?             @                     	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                      	          hff�?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @                                   �?8$�s���?�            `t@                                  @^@`'�J�?!            �I@                                  Pb@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                    �C@                                  �Z@X�)�O�?�            0q@        ������������������������       �        	             2@               T                   �z@���?�            p@               #       
             �?�X�<ݺ?�            �o@        !       "                   �r@ȵHPS!�?             :@       ������������������������       �                     7@        ������������������������       �                     @        $       C       	          ����?���=��?�            @l@       %       B                    �?@4և���?V            �_@       &       7                   @_@ �Cc}�?;             U@       '       6                   �[@�1�`jg�?'            �K@       (       1                    �? �Cc}�?             <@       )       *                    _@�����?             5@        ������������������������       �                     @        +       ,                   �Y@      �?             0@       ������������������������       �        	             $@        -       .                    @K@�q�q�?             @        ������������������������       �                     @        /       0                     Q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        2       3                   @^@؇���X�?             @        ������������������������       �                     @        4       5                   �Y@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        8       =                    `@V�a�� �?             =@        9       :                    @G@z�G�z�?             @        ������������������������       �                      @        ;       <                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        >       A                    b@�8��8��?             8@        ?       @                   �m@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     E@        D       E                    @J@p���?=             Y@        ������������������������       �                     D@        F       Q                    c@(;L]n�?'             N@       G       H       	             @0�)AU��?%            �L@       ������������������������       �                    �B@        I       P                   @^@P���Q�?             4@       J       K                    �?�����H�?             "@        ������������������������       �                     @        L       M                   �[@r�q��?             @        ������������������������       �                      @        N       O                     M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        R       S                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        U       V                   �X@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        X       o                    a@����+�?i            `d@        Y       h                   �r@�J�4�?0            �R@       Z       [                   @\@t�U����?*            �P@        ������������������������       �                     ;@        \       a                     P@z�G�z�?             D@       ]       `                   �`@ȵHPS!�?             :@       ^       _                    �?�θ�?	             *@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     *@        b       c                    �?X�Cc�?	             ,@        ������������������������       �                      @        d       e                   `c@      �?             (@       ������������������������       �                     @        f       g                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        i       n                     N@      �?              @       j       m       	          ����?�q�q�?             @       k       l                   `c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        p       {                    �?~�4_�g�?9             V@        q       z       	             @z�G�z�?             4@       r       u                   �a@�����H�?             2@        s       t                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        v       y       	          ����?@4և���?
             ,@        w       x                    @L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        |       }       
             �?      �?+             Q@        ������������������������       �                     $@        ~       �                   �`@�f7�z�?%             M@              �                    �?     ��?             @@       �       �                   �a@�θ�?             :@        ������������������������       �                      @        �       �       	          ���@r�q��?             8@       �       �                    �?�C��2(�?             6@        ������������������������       �                     @        �       �                    X@�t����?             1@        ������������������������       �                     �?        �       �                    @L@      �?
             0@       ������������������������       �                     "@        �       �       	          ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    @O@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?$�q-�?             :@       �       �                   Pr@`2U0*��?             9@       ������������������������       �                     8@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?>A�F<�?�            �w@       �       �                   @E@X��Oԣ�?�            `s@        �       �                   �]@���Q��?             4@        �       �                   @\@      �?             @       �       �                    [@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          `ff�?     ��?             0@        �       �       	          433�?r�q��?             @       ������������������������       �                     @        �       �                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�5�s��?�             r@        �       �                    �?b�h�d.�?,            �Q@        �       �                   �i@�G�z��?             4@        �       �                    `@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   ``@�q�q�?
             .@        �       �                   �[@����X�?             @        ������������������������       �                     �?        �       �                   �]@r�q��?             @        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    Z@ "��u�?             I@        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?`�q�0ܴ?            �G@       �       �                    b@�X�<ݺ?             B@       �       �                    ]@г�wY;�?             A@        �       �                   �[@      �?              @       ������������������������       �                     @        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �       �                     J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �t@P���Q�?�            �k@       �       �                    �?�6l�?�            `j@       �       �                   0h@ �.�?Ƞ?K             ^@       �       �                    �? 4^��?J            �]@        ������������������������       �                     E@        �       �                    @L@�e���@�?2            @S@       ������������������������       �        *             P@        �       �                   �_@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        �       �                     I@0�>���?:            �V@        �       �                    �?�*/�8V�?            �G@        �       �                   �d@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @[@Du9iH��?            �E@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        ������������������������       �                      F@        �       �                   �c@X�<ݚ�?             "@        �       �       	          ����?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   Pd@      �?)            �Q@       �       �                   �[@�^���U�?"            �L@        ������������������������       �                     @        �       �                    �?r�z-��?             �J@       �       �                    �?d}h���?             E@        ������������������������       �                     �?        �       �                   �`@��P���?            �D@       �       �                   �c@�G�z��?             4@       �       �                   ps@     ��?             0@       �       �                   �^@X�Cc�?	             ,@       �       �                    �?      �?             $@       �       �                     P@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             5@        �       �                    �?"pc�
�?             &@       ������������������������       �                     @        �       �                   �_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �T8q���?��cG��?�dn��i�?�f�P���?QFo�Z�?6��T��?����X�?^N��)x�?              �?|a���?�rO#,��?      �?        �;�;�?'vb'vb�?F]t�E�?]t�E�?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�q�q�?9��8���?      �?                      �?n�
�E�?P�T�;�?�?�������?UUUUUU�?�������?              �?      �?                      �?���ʭ?#�5�_#�?              �? ���?����?�q�q�?��8��8�?�؉�؉�?��N��N�?              �?      �?        Ź�Q��?d�:Fq�?�$I�$I�?n۶m۶�?۶m۶m�?%I�$I��?�־a�?A��)A�?۶m۶m�?%I�$I��?�a�a�?=��<���?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?a���{�?��{a�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?{�G�z�?\���(\�?              �?�?�������?p�}��?��Gp�?              �?�������?ffffff�?�q�q�?�q�q�?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?      �?                      �?[�o�W�?t�>H��?{�G�z�?�z�G��?g��1��?���-�?              �?�������?�������?�؉�؉�?��N��N�?�؉�؉�?ى�؉��?      �?                      �?              �?�m۶m��?%I�$I��?      �?              �?      �?              �?333333�?�������?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?              �?/�袋.�?��.���?�������?�������?�q�q�?�q�q�?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?      �?      �?      �?        a���{�?O#,�4��?      �?      �?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?]t�E�?F]t�E�?      �?        <<<<<<�?�?              �?      �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?{�G�z�?���Q��?              �?      �?              �?        ������?Cy�5��?c�1�c�?�s�9�?�������?333333�?      �?      �?      �?      �?      �?                      �?      �?              �?      �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?�d�&Jv�?��DɮM�?;��:���?_�_��?�������?�������?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �G�z�?���Q��?UUUUUU�?UUUUUU�?      �?                      �?��F}g��?W�+�ɥ?��8��8�?�q�q�?�?�?      �?      �?      �?              �?      �?      �?                      �?      �?              �?      �?      �?                      �?      �?        ffffff�?�������?�۩<:��?_Fb5\��?wwwwww�?�?�(��(��?�5�5�?      �?        qV~B���?�cj`?      �?        �؉�؉�?;�;��?              �?      �?                      �?��=��=�?�!�!�?r1����?m�w6�;�?      �?      �?              �?      �?        qG�w��?w�qGܱ?      �?      �?      �?                      �?      �?              �?        r�q��?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?:��,���?c:��,��?      �?        �琚`��?����!�?۶m۶m�?I�$I�$�?              �?�����?������?�������?�������?      �?      �?%I�$I��?�m۶m��?      �?      �?r�q��?�q�q�?      �?                      �?              �?      �?                      �?              �?              �?/�袋.�?F]t�E�?      �?              �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJKcChG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�G         �       	          033�?N�[7���?Y           ��@              +                   `^@N��y��?P           �@                      
             �?������?U             `@                                  �?h�˹�?5             S@                                 �]@�3Ea�$�?              G@                                  �?؇���X�?             E@                                   �K@z�G�z�?
             .@        ������������������������       �                     @        	       
                   �X@      �?              @        ������������������������       �                     @        ������������������������       �                     @                                  �Y@�����H�?             ;@        ������������������������       �        	             *@                      
             �?d}h���?             ,@        ������������������������       �                     �?                                   l@�θ�?
             *@       ������������������������       �                     @                      	          ����?      �?             @        ������������������������       �                     @        ������������������������       �                     @                                   �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     >@               $                   �S@�iʫ{�?             �J@                                  �]@��
ц��?             *@                                  �[@����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                   �?r�q��?             @        ������������������������       �                     �?                #                    �?z�G�z�?             @       !       "                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        %       &                    �?P���Q�?             D@       ������������������������       �                    �@@        '       (                   �p@����X�?             @       ������������������������       �                     @        )       *                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ,       ]                    �?     n�?�             x@        -       R                    �?�������?U             ^@       .       =       
             �?�"���r�?D            �X@        /       2                   �_@p9W��S�?             C@        0       1       	          ����?�X�<ݺ?             2@       ������������������������       �        
             1@        ������������������������       �                     �?        3       :                   �a@      �?             4@       4       5                    �?�	j*D�?
             *@        ������������������������       �                     @        6       9                    q@      �?              @       7       8       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ;       <                   �t@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        >       A                   �b@��6}��?)            �N@        ?       @                    �?Pa�	�?            �@@        ������������������������       �                     �?        ������������������������       �                     @@        B       I                    �I@���>4��?             <@        C       D                   �c@����X�?             ,@        ������������������������       �                     @        E       F                   pf@�C��2(�?	             &@       ������������������������       �                      @        G       H                    @E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        J       O                    �?d}h���?             ,@        K       L                   @d@      �?             @        ������������������������       �                     �?        M       N                   �_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        P       Q                   f@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        S       X                   pa@����X�?             5@        T       U                   a@����X�?             @        ������������������������       �                     @        V       W                   @[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        Y       Z                   0j@@4և���?             ,@       ������������������������       �                     "@        [       \                    ]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       w                    @L@���L:�?�            �p@       _       h       
             �?��S�ۿ?�            @j@        `       a                    �?
;&����?             7@        ������������������������       �                      @        b       c                    �C@������?             .@        ������������������������       �                     @        d       g       	          @33�?���|���?             &@       e       f                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        i       t                   h@Pհ�*�?v            `g@       j       m                    I@�����?t             g@        k       l                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        n       o                    �? Y@��?p            �f@       ������������������������       �        @            �X@        p       q                    �? �)���?0            @T@        ������������������������       �                     8@        r       s                   @[@0�)AU��?"            �L@        ������������������������       �                     �?        ������������������������       �        !             L@        u       v                    d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        x       �       
             �?�E��ӭ�?              K@        y       |                    �?ҳ�wY;�?	             1@        z       {                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        }       �                    �?����X�?             ,@       ~                           c@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?������?            �B@        �       �                    �?d}h���?             ,@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   0c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �L@ףp=
�?             $@        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   pa@�nkK�?             7@        ������������������������       �                     $@        �       �                    �?$�q-�?             *@       ������������������������       �                     $@        �       �       	          @33�?�q�q�?             @       �       �                   0d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �             
             �?_H���?	           Py@       �       �                    �?ZD�ɴ�?�            `u@        �       �                    �?��7��?$            �N@       �       �       	             �?����e��?            �@@       �       �                    �H@���N8�?             5@        ������������������������       �                      @        �       �       	             �?�S����?             3@        �       �                   �o@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                   Xr@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �_@�q�q�?             (@        �       �                    b@���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?؇���X�?             @        ������������������������       �                     �?        �       �                    �E@r�q��?             @        ������������������������       �                     @        �       �       	          `ff@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����? �Cc}�?             <@        ������������������������       �                     &@        �       �       	          ����?@�0�!��?
             1@        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        �       �                   `b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@4և���?             ,@       �       �                   Pj@؇���X�?             @        ������������������������       �                     @        �       �                    d@      �?             @       �       �                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �                         �z@��L��?�            �q@       �       �                    �? ���g=�?�            @q@       �       �                   �e@�:���ΰ?�            �i@       �       �                   �V@�)f5��?�            �i@        ������������������������       �                     �?        �       �                    �?0���{�?�            �i@       �       �                    �?@�z�G�?f             d@        �       �                   ``@XB���?             =@       ������������������������       �        
             3@        �       �                   pr@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                   �e@��"pK�?V            ``@        �       �                   @e@�g�y��?             ?@       ������������������������       �                     >@        ������������������������       �                     �?        ������������������������       �        ?             Y@        �       �                   �_@t��ճC�?              F@        �       �                   �^@և���X�?             @       �       �       
             �?z�G�z�?             @       ������������������������       �                     @        �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �B@        ������������������������       �                     �?        �                          e@X�Cc�?/            �Q@       �       �                    @F@�X����?-            �P@        �       �       	             @      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �       	             �?�c�Α�?&             M@        �       �                    �?r�q��?             >@       �       �       	             �?�q�q�?
             (@       �       �                    �?      �?             $@       �       �                   0r@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             2@        �       �       	          033�?��>4և�?             <@        �       �                   `@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @L@���!pc�?             6@        �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                   `a@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �             	          ���@z�G�z�?             .@       �       �                    �?և���X�?             @        ������������������������       �                      @        �                           �?���Q��?             @       �       �       	             @      �?             @        �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                ``@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @                                 �?�G��l��?+            �O@                                �F@6YE�t�?            �@@        	      
                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                �_@ףp=
�?             >@        ������������������������       �        
             .@                                 �?z�G�z�?             .@        ������������������������       �                     @                                 �?�z�G��?             $@                                �]@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                @b@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �M@r�q��?             >@                                �L@ �q�q�?             8@       ������������������������       �                     4@                                �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                �p@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �t�b��     h�h)h,K ��h.��R�(KMKK��hb�B�  �3��3��?f�f��?Q]Eu��?]Eu�U�?���-iK�?��-iK��?�5��P�?^Cy�5�?��,d!�?����7��?�$I�$I�?۶m۶m�?�������?�������?              �?      �?      �?      �?                      �?�q�q�?�q�q�?              �?۶m۶m�?I�$I�$�?              �?�؉�؉�?ى�؉��?              �?      �?      �?              �?      �?              �?      �?              �?      �?                      �?
�[���?�琚`��?�؉�؉�?�;�;�?�m۶m��?�$I�$I�?              �?      �?        UUUUUU�?�������?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?ffffff�?�������?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?             ��?      �?�������?�������?ogH���?"1ogH��?l(�����?�k(����?�q�q�?��8��8�?              �?      �?              �?      �?vb'vb'�?;�;��?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        �!XG��?;ڼOq��?|���?|���?              �?      �?        n۶m۶�?I�$I�$�?�m۶m��?�$I�$I�?              �?]t�E�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?I�$I�$�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?        �$I�$I�?�m۶m��?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?        �$I�$I�?n۶m۶�?              �?�������?�������?      �?                      �?|��|�?|���?�������?�?Y�B��?�Mozӛ�?      �?        �?wwwwww�?              �?F]t�E�?]t�E]�?�q�q�?9��8���?      �?                      �?      �?        }�ٓ|�?n�ʄm�?zӛ����?d!Y�B�?      �?      �?      �?                      �?(}�'}��?l�l�v?      �?        X�<ݚ�?�����H�?      �?        ��Gp�?p�}��?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�q�q�?r�q��?�������?�������?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?              �?      �?                      �?��g�`��?к����?I�$I�$�?۶m۶m�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?      �?                      �?      �?        �Mozӛ�?d!Y�B�?      �?        �؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �g�����?�D��?R[Im%��?+������?�y��!�?&C��6��?e�M6�d�?6�d�M6�?�a�a�?��y��y�?              �?(������?^Cy�5�?      �?      �?      �?        �������?333333�?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?%I�$I��?              �?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�$I�$I�?n۶m۶�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?      �?      �?                      �?              �?              �?�\���?����?ہ�v`��?��(�3J�?�H%�e�?�~�����?��߁��?��;�?      �?        �?777777�?�������?�������?�{a���?GX�i���?              �?�������?�������?              �?      �?        qBJ�eD?{k�4w��?�B!��?��{���?              �?      �?                      �?t�E]t�?�E]t��?۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?      �?                      �?      �?                      �?      �?        �m۶m��?%I�$I��?]t�E]�?�E]t��?      �?      �?      �?                      �?�{a���?5�rO#,�?UUUUUU�?�������?�������?�������?      �?      �?UUUUUU�?�������?              �?      �?              �?                      �?              �?I�$I�$�?۶m۶m�?�������?UUUUUU�?      �?                      �?t�E]t�?F]t�E�?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?        �������?�������?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?      �?        333333�?�������?              �?      �?        ��y��y�?1�0��?e�M6�d�?'�l��&�?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?�������?�������?              �?333333�?ffffff�?      �?      �?              �?      �?        UUUUUU�?�������?      �?                      �?�������?UUUUUU�?�������?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJN]{hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@C         z                   �`@��J�0�?B           ��@               =       	             �?�1�C��?           `|@                                  �S@�0u��A�?u            �f@                      
             �?R�(CW�?3            �T@                     	          033�?��GEI_�?'            �N@                                  @L@h�����?$             L@                                   @K@$�q-�?             :@       ������������������������       �                     5@        	       
                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     >@                      
             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                   �?և���X�?             5@                                 �c@      �?	             2@                                 @_@���Q��?             .@                                  �?�q�q�?             "@                                  \@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               ,                    �?և���X�?B            �X@              #                    �?.��<�?/            �P@                                   @Y@����X�?             5@                                  �k@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        !       "       
             �?�r����?
             .@       ������������������������       �                     *@        ������������������������       �                      @        $       +                   �~@�nkK�?              G@       %       *       
             �?����?�?            �F@        &       )       	          ����?�q�q�?             @       '       (                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     E@        ������������������������       �                     �?        -       .                    [@�n`���?             ?@        ������������������������       �                     �?        /       8       	          ����?r�q��?             >@       0       5                   `q@H%u��?             9@       1       4                    �?���7�?             6@        2       3                    �J@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     (@        6       7                   @_@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        9       <       	          ����?���Q��?             @       :       ;                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        >       ?                   �Q@DS���|�?�             q@        ������������������������       �                      @        @       U                    @M@�?�0�!�?�             q@       A       L       	          ����?����=O�?T             b@        B       K                    @�?�'�@�?             C@       C       F                    �?������?            �B@        D       E                   �e@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        G       H                    �?      �?             @@       ������������������������       �                     >@        I       J                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        M       T       	          ����?���1��??            �Z@        N       S                    \@г�wY;�?             A@        O       R                   m@؇���X�?             @        P       Q                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        ������������������������       �        *            @R@        V       _                    �M@�'F����?I            �_@        W       ^                    �?      �?
             4@       X       Y                   �_@�q�q�?             .@        ������������������������       �                      @        Z       [       
             �?�θ�?             *@        ������������������������       �                      @        \       ]                   �]@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        `       w                    �R@��hq��??            �Z@       a       n                   p`@�b�E�V�?<            �Y@        b       k                    �?@�0�!��?             A@       c       d                   �Y@     ��?             0@        ������������������������       �                      @        e       f                   �q@d}h���?             ,@       ������������������������       �                      @        g       h                   �_@      �?             @        ������������������������       �                      @        i       j                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        l       m                    �?�X�<ݺ?	             2@       ������������������������       �                     1@        ������������������������       �                     �?        o       p                   pb@��.N"Ҭ?&            @Q@       ������������������������       �                    �G@        q       r                    `P@�C��2(�?             6@       ������������������������       �                     *@        s       t                   �N@�<ݚ�?             "@        ������������������������       �                     �?        u       v                    �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        x       y       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        {       �       
             �?n���?/            }@        |       �                    �?�E�Y��?x            �g@       }       �                    �?؇���X�?C            @Z@        ~       �                   �a@      �?             8@              �                    �?���Q��?             .@       �       �                    �?      �?             (@        ������������������������       �                     @        �       �                   �a@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�����H�?5            @T@        �       �                    �?�r����?             >@       �       �                   �e@��s����?             5@       �       �       
             �?�KM�]�?             3@        ������������������������       �                     �?        �       �                   �`@�����H�?             2@       �       �                   xr@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    \@`�H�/��?            �I@        �       �                   �m@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?���.�6�?             G@        ������������������������       �                     (@        �       �                   0c@l��\��?             A@       ������������������������       �                     ;@        �       �                     M@և���X�?             @        ������������������������       �                      @        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �P@`m:*G��?5            �U@       �       �                    �?�ҿf���?3            �T@        �       �       	          033@l��
I��?             ;@       �       �                   �q@�GN�z�?             6@       �       �       	          ����?      �?             0@        �       �                    �N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@        �       �                   `]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?���>4��?"             L@        ������������������������       �                     @        �       �       	          ����?X�Emq�?!            �J@        �       �                     G@@�0�!��?
             1@        ������������������������       �                     @        ������������������������       �                     ,@        �       �                    �I@X�<ݚ�?             B@       �       �                   �f@��Q��?             4@       �       �       	             @������?             1@       �       �                   �`@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   Po@     ��?
             0@       �       �                   �l@�8��8��?             (@       ������������������������       �                     @        �       �                    n@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �p@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?R��N�?�            q@        �       �                   a@F�����?            �F@        ������������������������       �                     @        �       �                    �?v�2t5�?            �D@        ������������������������       �        	             *@        �       �                    @G@��>4և�?             <@        �       �                    �?�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pb@�<ݚ�?             2@        �       �                    �O@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �K@8�Z$���?             *@        �       �                   �n@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   @E@h�˹�?�            �l@        �       �                   @Z@������?             1@        �       �       	          ���Ὸ��Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �b@�8��8��?
             (@        ������������������������       �                     @        �       �       	          433�?z�G�z�?             @       ������������������������       �                     @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                          �?`[ү��?�            `j@       �       �                    �?��I�~R�?�            �h@        �       �                   pf@R���Q�?             D@       �       �                   �_@������?            �B@        �       �                   Po@������?             1@       �       �                    �?�r����?
             .@       �       �       	          ����?8�Z$���?	             *@       �       �                   pl@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                   pe@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     4@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �^@�#��g1�?j            �c@        ������������������������       �        $             K@        �                          _@ f^8���?F            �Y@        �                           �?���Q��?             @       �       �                   �l@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                 �?@uvI��?C            �X@       ������������������������       �        $            �K@                                pa@ qP��B�?            �E@       ������������������������       �                     <@                                �r@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        	      
      	          `ff�?X�Cc�?	             ,@        ������������������������       �                      @                                �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  �̓"��?�6�n��?H@ͮY�?�L�)�?�������?�������?KԮD�J�?�JԮD��?;ڼOqɰ?�d����?�$I�$I�?�m۶m��?;�;��?�؉�؉�?              �?�������?333333�?      �?                      �?              �?�������?333333�?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?                      �?              �?�$I�$I�?۶m۶m�?IT�n��?o�Wc"=�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?�?�������?              �?      �?        �Mozӛ�?d!Y�B�?��I��I�?l�l��?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?�c�1��?�9�s��?      �?        UUUUUU�?�������?���Q��?)\���(�?F]t�E�?�.�袋�?�������?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?�uy)�?I�ܺ�?      �?        xxxxxx�?�������?��RA�/�?U��K��?y�5���?������?к����?��g�`��?333333�?�������?              �?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        �+J�#�?�S�rp��?�?�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?              �?              �?
�B�P(�?�^�����?      �?      �?UUUUUU�?UUUUUU�?              �?ى�؉��?�؉�؉�?              �?]t�E�?F]t�E�?              �?      �?                      �?�Ե��?bEi|d�?��,�?�jch���?�������?ZZZZZZ�?      �?      �?      �?        ۶m۶m�?I�$I�$�?              �?      �?      �?              �?      �?      �?      �?                      �?�q�q�?��8��8�?              �?      �?        ہ�v`��?�3J���?              �?F]t�E�?]t�E�?              �?�q�q�?9��8���?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?��FX��?�4�rO#�?�d�h��?�M�˘��?�$I�$I�?۶m۶m�?      �?      �?�������?333333�?      �?      �?      �?              �?      �?      �?                      �?              �?              �?�q�q�?�q�q�?�?�������?�a�a�?z��y���?(�����?�k(���?              �?�q�q�?�q�q�?      �?      �?              �?      �?              �?      �?              �?      �?              �?                      �?�?�������?�������?333333�?      �?                      �?Y�B��?���7���?              �?�������?------�?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?                      �?0�����?�/����?S��rY�?Y1P�M�?Lh/����?h/�����?�袋.��?]t�E�?      �?      �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?              �?      �?        n۶m۶�?I�$I�$�?      �?        �}�	��?5�x+��?�������?ZZZZZZ�?      �?                      �?r�q��?�q�q�?ffffff�?�������?�?xxxxxx�?F]t�E�?]t�E]�?      �?                      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?      �?              �?      �?                      �?{��z���?J�J��?�>�>��?؂-؂-�?      �?        ��+Q��?�ڕ�]��?      �?        I�$I�$�?۶m۶m�?ffffff�?333333�?              �?      �?        �q�q�?9��8���?�������?333333�?              �?      �?        ;�;��?;�;��?�������?333333�?      �?                      �?              �?^Cy�5�?�5��P�?�?xxxxxx�?333333�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?      �?              �?      �?        4�Syt��?_Fb5\��?�Y���?\e
�d�?333333�?333333�?��g�`��?к����?xxxxxx�?�?�������?�?;�;��?;�;��?]t�E�?F]t�E�?      �?                      �?      �?      �?              �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?>"'wc�?A����?      �?        H%�e�?��VCӝ?333333�?�������?      �?      �?      �?                      �?      �?        �Cc}h��?9/���?      �?        ��}A�?�}A_З?      �?        �������?�?      �?                      �?%I�$I��?�m۶m��?      �?        UUUUUU�?�������?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�|�7hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@G         z                   a@z�ГPo�?T           ��@               ;                    �?�����?&           �|@               &       
             �?�s���?s             f@              !                   �r@
��^���?<            @W@                                 `\@�~6�]�?6            @U@                                   �?��?^�k�?            �A@                                   �?��S�ۿ?
             .@       ������������������������       �                     $@        	              	          @33�?z�G�z�?             @       
                          �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@                                   �?�w��#��?             I@                                   �?z�G�z�?             $@                                   �J@      �?             @        ������������������������       �                     �?                                  @k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                  @L@R���Q�?             D@                      	          `ff�?���Q��?
             4@        ������������������������       �                     @                                   �?�n_Y�K�?             *@        ������������������������       �                      @        ������������������������       �                     @                                    @F@P���Q�?             4@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        "       #                    @G@      �?              @        ������������������������       �                      @        $       %       	          ���@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        '       6       	          ����?d}h���?7             U@       (       1                    �?�L#���?-            �P@        )       0                   �_@@�0�!��?             1@       *       +                    �?�q�q�?             "@        ������������������������       �                      @        ,       -                   `[@և���X�?             @        ������������������������       �                     @        .       /                    �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        2       3                   `c@p���?             I@       ������������������������       �                     G@        4       5                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        7       8                   �e@@�0�!��?
             1@       ������������������������       �                     *@        9       :       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        <       c                   P`@���J�?�            �q@        =       \                    �?��j���?J            �[@       >       Y                   0r@�:nR&y�?B            �W@       ?       V                     R@������?:            �T@       @       A                    �?x�G�z�?8             T@        ������������������������       �                     4@        B       K                   �_@P���Q�?(             N@       C       D                    @L@ ���J��?            �C@       ������������������������       �                     5@        E       F       	          033�?�X�<ݺ?             2@       ������������������������       �                     $@        G       H       
             �?      �?              @        ������������������������       �                     @        I       J       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        L       U                    �?�����?             5@       M       T       	          ����?      �?             0@        N       S                   �[@���Q��?             @       O       P                    `@�q�q�?             @        ������������������������       �                     �?        Q       R                   �Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        W       X                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Z       [                   �r@�θ�?             *@        ������������������������       �                     @        ������������������������       �                     $@        ]       b                   �]@      �?             0@       ^       a                     P@�q�q�?             "@       _       `                     F@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        d       q       
             �?蹱f
@�?i            �e@       e       p                   �b@�Fǌ��?^            �c@       f       g                   Pl@ _�@�Y�?G             ]@       ������������������������       �        '            �P@        h       m                   �b@@9G��?             �H@       i       l       	             �? qP��B�?            �E@        j       k                   `m@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        n       o                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     E@        r       y                   �^@��S���?             .@       s       x                    �?�n_Y�K�?	             *@       t       w       	             �?z�G�z�?             $@        u       v                   @\@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        {       �                    �K@T!y<�-�?.           �|@       |       �                    �?���@��?�            �r@        }       �                   �a@և���X�?E            @Z@        ~       �                    �?$��m��?             :@              �                   �\@�r����?             .@        ������������������������       �                     @        �       �       
             �?�<ݚ�?             "@        �       �                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?���|���?             &@       �       �                   �\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    f@H���I�?2            �S@       �       �       	          ����?|�U&k�?.            �R@       �       �                    �?և���X�?            �H@        ������������������������       �                     @        �       �                    �?���|���?             F@       �       �                    �?      �?             @@       �       �                   @_@�n_Y�K�?             :@        �       �                    �B@���|���?             &@        ������������������������       �                      @        �       �                   �[@�<ݚ�?             "@        �       �                   �g@���Q��?             @        ������������������������       �                      @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�G�z�?             .@       �       �       
             �?d}h���?             ,@        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?HP�s��?             9@        �       �       	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?���7�?             6@       �       �       
             �?ףp=
�?             $@        ������������������������       �                      @        �       �                    n@      �?              @        �       �       	             @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        �       �                    �?�8��8��?�             h@        �       �                    �?0�,���?)            �P@       �       �                   @a@ ������?&            �O@       ������������������������       �                     G@        �       �                     H@�IєX�?             1@       ������������������������       �                     $@        �       �                   p@؇���X�?             @        ������������������������       �                     @        �       �       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �_@      �?             @        ������������������������       �                      @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �g@Tb.��?W            @_@       �       �       
             �?�חF�P�?V             _@        �       �                   ``@��X��?             <@       �       �                    �?��S���?             .@        ������������������������       �                     @        �       �                   @Z@�z�G��?             $@        ������������������������       �                     �?        �       �                     G@�<ݚ�?             "@       �       �                     B@���Q��?             @        ������������������������       �                      @        �       �                   @_@�q�q�?             @       �       �                    �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   pr@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �       	          ���@�q�q�?A             X@       ������������������������       �        @            �W@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��Q�e�?i             d@        �       �                    �?.�	F�9�?4            @T@       �       �                    �?��U/��?$            �L@        �       �                   `a@��2(&�?             6@        ������������������������       �                      @        �       �                   �v@P���Q�?             4@       ������������������������       �                     .@        �       �       	          ���@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?���Q��?            �A@        �       �                   g@d}h���?	             ,@        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          @33�?�C��2(�?             &@        �       �                   �b@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   c@؇���X�?             5@       �       �                   �p@�IєX�?             1@       ������������������������       �                     (@        �       �                   �_@z�G�z�?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     8@        �       
                  �b@v�_���?5            �S@        �       �       	          @33�?X�<ݚ�?             B@        �       �                   �`@ףp=
�?             $@        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                 m@R�}e�.�?             :@                                `Z@      �?             (@        ������������������������       �                     @                                �a@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?              	                   �?@4և���?	             ,@                    
             �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@                                 @�T|n�q�?            �E@                   	             @ףp=
�?             >@                               �`@@4և���?             <@        ������������������������       �                     $@                                hs@�����H�?             2@       ������������������������       �        
             ,@                                  P@      �?             @        ������������������������       �                      @        ������������������������       �                      @                    	             @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                �e@�	j*D�?             *@                   	          033�?"pc�
�?             &@                                 �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  1�i�M��?��<Y �? ��:��?8�Hq�?�F($�?Cr����?��~���?X`��?�?999999�?�A�A�?_�_��?�?�������?              �?�������?�������?      �?      �?      �?                      �?              �?              �?��(\���?��Q��?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?�������?333333�?              �?;�;��?ى�؉��?      �?                      �?�������?ffffff�?      �?      �?      �?                      �?              �?      �?      �?              �?�������?UUUUUU�?      �?                      �?I�$I�$�?۶m۶m�?��@���?g��1��?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?              �?        \���(\�?{�G�z�?      �?              �?      �?              �?      �?        �������?ZZZZZZ�?              �?      �?      �?      �?                      �?��RO�o�?A�6�?�9	ą��?����^�?�-q��ܲ?Fڱa��?������?p>�cp�?333333�?�������?              �?�������?ffffff�?�A�A�?��-��-�?              �?�q�q�?��8��8�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�a�a�?=��<���?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?              �?      �?      �?      �?                      �?�؉�؉�?ى�؉��?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?        \
�IƢ�?Z/`��U�?�3���?1���M��?�{a���?#,�4�r�?              �?9/���?������?�}A_З?��}A�?      �?      �?      �?                      �?              �?UUUUUU�?�������?      �?                      �?              �?�������?�?ى�؉��?;�;��?�������?�������?      �?      �?              �?      �?                      �?      �?              �?        �0�����?��=^�?H�8��?q5���?۶m۶m�?�$I�$I�?�N��N��?vb'vb'�?�������?�?      �?        9��8���?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?        F]t�E�?]t�E]�?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?      �?                      �?^-n����?Q�Ȟ���?E>�S��?�`�|��?۶m۶m�?�$I�$I�?      �?        F]t�E�?]t�E]�?      �?      �?;�;��?ى�؉��?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?I�$I�$�?۶m۶m�?              �?      �?              �?                      �?              �?{�G�z�?q=
ףp�?UUUUUU�?UUUUUU�?              �?      �?        F]t�E�?�.�袋�?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �����*�?�������?Ez�rv�?g��1��?��}��}�?AA�?      �?        �?�?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?      �?              �?      �?              �?      �?        9��v���?/�$��?�Zk����?��RJ)��?%I�$I��?n۶m۶�?�?�������?      �?        333333�?ffffff�?      �?        �q�q�?9��8���?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?;�;��?�؉�؉�?              �?      �?        �������?UUUUUU�?      �?                      �?              �?�������?333333�?~X�<��?�����H�?g1��t�?Lg1��t�?t�E]t�?��.���?      �?        �������?ffffff�?              �?�������?�������?      �?                      �?�������?333333�?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?]t�E�?F]t�E�?�������?�������?              �?      �?              �?        �$I�$I�?۶m۶m�?�?�?              �?�������?�������?              �?      �?      �?              �?      �?              �?      �?              �?      �?                      �? *�3�?���M���?�q�q�?r�q��?�������?�������?      �?        �������?�������?      �?                      �?�;�;�?'vb'vb�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?                      �?�$I�$I�?n۶m۶�?�������?�������?              �?      �?                      �?���)k��?6eMYS��?�������?�������?n۶m۶�?�$I�$I�?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?              �?      �?              �?      �?        vb'vb'�?;�;��?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJsO�'hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         n                   p`@�7i���?5           ��@               ;                    �?���ě)�?�            @y@               *       
             �?� �	��?_            �b@                                  �?��܂O�?8            �V@                                   �?d}h���?             ,@                                 `j@�8��8��?             (@        ������������������������       �                      @               	                   �a@      �?             @        ������������������������       �                      @        
              	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @               !                     Q@�C��2(�?0            @S@                                  �? =[y��?)             Q@                                 �k@�O4R���?             �J@       ������������������������       �                     @@                                  �k@���N8�?             5@                                   �?r�q��?             @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@                                    a@�r����?	             .@                     
             �?����X�?             @        ������������������������       �                     �?                                  `X@r�q��?             @                                   @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        "       )                    @R@X�<ݚ�?             "@       #       (       	          ����?�q�q�?             @       $       %                    b@�q�q�?             @        ������������������������       �                     �?        &       '                   Pf@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        +       :                    @F�4�Dj�?'            �M@       ,       3                    �?؇���X�?$             L@       -       2                    �?dP-���?            �G@        .       1                   �_@������?             .@        /       0                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @@        4       9                    �?X�<ݚ�?             "@       5       8                    �?����X�?             @       6       7       	          @33�?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        <       i                   �e@R�xE��?�            �o@       =       f                    @أ����?�            �n@       >       _       
             �?���X=P�?�            �n@       ?       @                   Pe@�j�-��?�            `l@        ������������������������       �        0            @S@        A       L                    `@���Lͩ�?X            �b@        B       K                    �?r�q��?             E@       C       D                   8p@      �?             D@       ������������������������       �                     5@        E       J                   �_@�d�����?             3@       F       G                    �?      �?
             0@       ������������������������       �                     (@        H       I                    Z@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        M       N                   �e@��Wv��?>             [@        ������������������������       �                     @        O       ^                    �R@��FM ò?=            @Z@       P       U                    @H@p� V�?<            �Y@        Q       R                   Pl@��S�ۿ?
             .@        ������������������������       �                     @        S       T       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        V       ]                    �L@�|���?2             V@        W       X                    @L@P�Lt�<�?             C@       ������������������������       �                     >@        Y       \                    Z@      �?              @        Z       [                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     I@        ������������������������       �                      @        `       a                    �?�E��ӭ�?             2@        ������������������������       �                     @        b       c                    �?�r����?	             .@       ������������������������       �                      @        d       e                     P@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        g       h                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        j       m       
             �?և���X�?             @       k       l                     L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        o       �                    �?��9��3�?>           �@        p       �                    �?4�3p1�?z            @i@       q       �                   �b@�`���?V            `b@       r       y                    [@d��0u��?4            �V@        s       t                    �?�z�G��?             $@        ������������������������       �                     @        u       v       
             �?      �?             @        ������������������������       �                      @        w       x                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        z       �                    �?�G�z�?/             T@        {       �                   0a@     ��?             @@       |       �                   �`@\X��t�?             7@       }       �                   hp@�ՙ/�?             5@       ~                          �[@���!pc�?             &@        ������������������������       �                     �?        �       �                    �F@z�G�z�?             $@        ������������������������       �                     �?        �       �                   �`@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                     "@        �       �       
             �?�8��8��?             H@       �       �                   �m@��Y��]�?            �D@        �       �                    �G@�}�+r��?
             3@        �       �                   �k@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     6@        �       �       	          ����?և���X�?             @        ������������������������       �                      @        �       �       	          033�?z�G�z�?             @        ������������������������       �                     @        �       �                   `W@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �e@�����?"            �L@       �       �                   �d@���Q��?            �F@       �       �                   �i@���!pc�?            �@@        �       �                    �O@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?PN��T'�?             ;@       �       �       	          `ff@HP�s��?             9@       ������������������������       �                     7@        ������������������������       �                      @        ������������������������       �                      @        �       �                   �u@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?�C��2(�?$            �K@        �       �                    a@      �?             (@        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?             @        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pa@ �#�Ѵ�?            �E@        �       �                    �M@���Q��?             @       �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     C@        �       �       
             �?:�&���?�            �s@        �       �                   �Q@ܐ҆��?<            @W@        ������������������������       �                     @        �       �                   �l@������?7            �U@        �       �                   �_@�z�G��?             D@       ������������������������       �                     0@        �       �                   `a@      �?             8@        �       �                    j@�q�q�?             (@        ������������������������       �                     @        �       �                   �`@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             (@        ������������������������       �                      @        �       �                   �d@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                   f@��C���?             �G@       �       �       
             �?�E��ӭ�?             B@        �       �                   �l@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `]@     ��?             @@        ������������������������       �                     @        �       �                    �H@R�}e�.�?             :@        ������������������������       �                     @        �       �                   �q@��Q��?             4@       �       �                   @e@      �?
             ,@       �       �                    �?���|���?	             &@       �       �                   `d@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �N@���Q��?             @       �       �                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   pm@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                   0h@���O�?�            `k@       �       �                    �?�~�y�C�?�            @k@        �       �                     L@�LQ�1	�?             7@       ������������������������       �                     0@        �       �                   @a@և���X�?             @       �       �       	          ����?���Q��?             @       �       �                   �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    @L@��ɉ�?t            `h@       �       �       	             @@��'��?`             d@       ������������������������       �        _            �c@        ������������������������       �                      @        �       �                   �O@�t����?             A@        ������������������������       �                      @        �       �                   �d@      �?             @@       �       �                    �L@�����?             5@        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    d@�}�+r��?             3@       ������������������������       �        
             0@        �       �       	          833�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �t�b��:     h�h)h,K ��h.��R�(KK�KK��hb�B�  }}}}}}�?AAAAAA�?��N̓�?^?[���?)\���(�?�Q����?�Q�Q�?�������?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?              �?      �?                      �?F]t�E�?]t�E�?�������?�������?�x+�R�?:�&oe�?              �?�a�a�?��y��y�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�������?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?�q�q�?r�q��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?��/���?�A�I��?۶m۶m�?�$I�$I�?�����F�?W�+�ɵ?wwwwww�?�?r�q��?�q�q�?      �?                      �?      �?              �?        r�q��?�q�q�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?��`0�?>������?�KA���?���h�?]�l8bڳ?�j򸳄�?{��U���?覤:��?              �?�K~��?�6�i�?UUUUUU�?�������?      �?      �?              �?y�5���?Cy�5��?      �?      �?              �?      �?      �?              �?      �?              �?              �?        {	�%���?�^B{	��?      �?        8�8��?��~���?��,�?����`�?�?�������?              �?      �?      �?      �?                      �?F]t�E�?��.���?(�����?���k(�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        r�q��?�q�q�?      �?        �?�������?              �?�$I�$I�?�m۶m��?      �?                      �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?E�D�D��?w�v�v��?B���be�?߈�N��?և���X�?����S�?wwwwww�?DDDDDD�?ffffff�?333333�?      �?              �?      �?      �?              �?      �?      �?                      �?�������?�������?      �?      �?!Y�B�?��Moz��?�<��<��?�a�a�?t�E]t�?F]t�E�?      �?        �������?�������?      �?        �q�q�?�q�q�?      �?                      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?������?8��18�?(�����?�5��P�?�������?�������?              �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?      �?                      �?Q^Cy��?^Cy�5�?333333�?�������?F]t�E�?t�E]t�?UUUUUU�?�������?              �?      �?        &���^B�?h/�����?q=
ףp�?{�G�z�?      �?                      �?              �?      �?      �?              �?      �?              �?        F]t�E�?]t�E�?      �?      �?�������?333333�?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�}A_Ч?�/����?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�A�A�?�o��o��?,��,�?��~���?              �?�/�I�?��֡�l�?ffffff�?333333�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        g���Q��?L� &W�?r�q��?�q�q�?      �?      �?              �?      �?              �?      �?              �?�;�;�?'vb'vb�?              �?ffffff�?�������?      �?      �?]t�E]�?F]t�E�?�������?UUUUUU�?      �?                      �?�������?333333�?      �?      �?              �?      �?              �?                      �?              �?/�袋.�?F]t�E�?              �?      �?        ��{���?vA�a�?��Ṱ�?4R1�:#�?��Moz��?Y�B��?      �?        �$I�$I�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ?�?��? �����?�l<��?r���p�?      �?                      �?<<<<<<�?�?              �?      �?      �?=��<���?�a�a�?      �?      �?      �?                      �?�5��P�?(�����?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ9whG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKۅ�h��B�6         |                   �b@��3����?=           ��@              A                    �?�Ǧ��?�           p�@                                  P@�E��
��?�            �s@                                   �?>A�F<�?/             S@                                  �b@`՟�G��?             ?@                                  �?�f7�z�?             =@                     	             �?�z�G��?             4@              	                   �Z@�<ݚ�?
             2@        ������������������������       �                      @        
                          @\@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                   X@�q�q�?             "@        ������������������������       �                      @                                    J@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �F@               4       	          pff�?6�iL�?�            �m@              1                     R@�T��8��?~             h@              ,       
             �?��C�/��?{            `g@                      	          ����?�q�����?"             I@                                  �?���B���?             :@        ������������������������       �                     @                                  �`@���}<S�?             7@       ������������������������       �                     *@                                   @E@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @                +                   �b@�q�q�?             8@       !       "                    l@�����?             5@        ������������������������       �                     $@        #       *                   �_@"pc�
�?             &@        $       '                    �?���Q��?             @        %       &                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        (       )                    X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        -       0                    �?��[����?Y             a@        .       /                    @H@�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �        L            �]@        2       3       	          ����?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        5       :                    �?�%^�?            �E@        6       9                   `c@z�G�z�?             $@       7       8                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ;       <       
             �?�C��2(�?            �@@       ������������������������       �                     =@        =       >                   `a@      �?             @        ������������������������       �                      @        ?       @                    @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        B       w                    �?6uH���?�            `s@       C       v                    �N@$]^z���?�             m@       D       i       	          ����?؇���X�?i             d@       E       F                    U@�θ�?9            �V@        ������������������������       �                      @        G       h                   �a@���*~�?8            @V@       H       a       
             �?:���u��?/            @S@       I       J                    �C@8�Z$���?'            @P@        ������������������������       �                      @        K       L                    @G@�k�'7��?$            �L@        ������������������������       �                     @        M       N                   �f@H�ՠ&��?"             K@        ������������������������       �        	             .@        O       P       	          hff�?:�&���?            �C@        ������������������������       �                     &@        Q       R                   @Z@      �?             <@        ������������������������       �                      @        S       T                   0j@���B���?             :@        ������������������������       �                     �?        U       Z                   r@�J�4�?             9@       V       Y                   �l@��S�ۿ?             .@        W       X                   a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        [       \                   �\@�z�G��?             $@        ������������������������       �                     @        ]       `                    �?և���X�?             @       ^       _                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        b       g                    �?      �?             (@        c       d       	          ����?���Q��?             @        ������������������������       �                     �?        e       f                   0n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             (@        j       o                    �?��?^�k�?0            �Q@        k       n       	          ���@      �?             @       l       m                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        p       u                   �T@����e��?-            �P@        q       r                   �`@r�q��?             @       ������������������������       �                     @        s       t       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        (             N@        ������������������������       �        (            �Q@        x       {                    \@ ���J��?+            �S@        y       z                   �Z@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        '             R@        }       ~                   �O@      �?�            �r@        ������������������������       �                     (@               �                    �?����?�            �q@        �       �       	            �?4���C�?-            �P@       �       �                   ``@�G��l��?             E@       �       �                    c@��X��?             <@        ������������������������       �                      @        �       �                   @f@R�}e�.�?             :@       �       �                    @K@�+e�X�?             9@       �       �                    �B@�r����?
             .@        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?$�q-�?             *@        ������������������������       �                      @        �       �                   �[@�C��2(�?             &@        �       �       
             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �r@���Q��?             $@       �       �                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?@4և���?
             ,@        �       �                    b@r�q��?             @       ������������������������       �                     @        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   @e@      �?             8@       ������������������������       �                     1@        �       �                   �e@؇���X�?             @        �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �f@�~i��?�            @k@       �       �                    �?8��?�A�?�             k@        �       �       	          ����?�}�+r��?-             S@       �       �       
             �?�:�]��?            �I@        �       �                    �E@և���X�?             @        ������������������������       �                      @        �       �                   �a@���Q��?             @       �       �                    �?      �?             @       �       �                    e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?`���i��?             F@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �C@        ������������������������       �                     9@        �       �                    ]@`	�<��?T            �a@        �       �                    �?�X����?             6@        �       �       	          hff�?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                     F@      �?             (@        ������������������������       �                     @        �       �                     J@      �?              @        ������������������������       �                     @        �       �                   `m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?�D�d@6�?G            �]@        �       �                   0g@�t����?             A@        ������������������������       �                     @        �       �                    �?z�G�z�?             >@       �       �       
             �?؇���X�?             <@        ������������������������       �                      @        �       �                    @C@z�G�z�?             4@        ������������������������       �                     �?        �       �                   �`@�S����?             3@       ������������������������       �                     $@        �       �                   @b@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   Pd@�D�e���?1            @U@        �       �                   �t@�C��2(�?             6@       �       �                    d@���N8�?             5@       ������������������������       �                     2@        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        "            �O@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  iL��/�?�Y=v��?�)���?kr�
%�?;�;��?��؉���?Cy�5��?������?�s�9��?�1�c��?a���{�?O#,�4��?333333�?ffffff�?�q�q�?9��8���?              �?�������?333333�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?              �?      �?              �?                      �?ylE�pR�?'u_[�?�­���?��H	9�?a�2a�?{��c5{�?���Q��?�p=
ף�?ى�؉��?��؉���?      �?        d!Y�B�?ӛ���7�?              �?�������?�������?      �?                      �?UUUUUU�?�������?=��<���?�a�a�?      �?        /�袋.�?F]t�E�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?                      �?�8R4��?������}?��8��8�?�q�q�?              �?      �?              �?        UUUUUU�?�������?              �?      �?        �}A_�?�}A_��?�������?�������?�q�q�?�q�q�?      �?                      �?              �?F]t�E�?]t�E�?              �?      �?      �?      �?              �?      �?      �?                      �?��RJ)��?k���Zk�?��{a�?�=�����?�$I�$I�?۶m۶m�?�؉�؉�?ى�؉��?      �?        ��MmjS�?���d%+�?qV~B���?dj`��?;�;��?;�;��?              �?Lg1��t�?-����b�?      �?        {	�%���?������?              �?�o��o��?�A�A�?              �?      �?      �?      �?        ى�؉��?��؉���?      �?        {�G�z�?�z�G��?�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?ffffff�?              �?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?              �?      �?�������?333333�?      �?              �?      �?      �?                      �?      �?                      �?�A�A�?_�_��?      �?      �?      �?      �?      �?                      �?              �?|���?�>����?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?              �?�A�A�?��-��-�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?s �
��?2~�ԓ��?'�l��&�?m��&�l�?1�0��?��y��y�?%I�$I��?n۶m۶�?      �?        �;�;�?'vb'vb�?���Q��?R���Q�?�?�������?      �?      �?      �?                      �?;�;��?�؉�؉�?              �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        ��w� z�?��A��.�?�nr7���?وlD6"�?�5��P�?(�����?}}}}}}�?�?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?      �?      �?      �?                      �?              �?      �?        F]t�E�?F]t�E�?�������?�������?              �?      �?              �?              �?        o����?E�)͋?�?�E]t��?]t�E]�?�������?�������?      �?                      �?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        }��|���?���й?�������?�������?              �?�������?�������?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?(������?^Cy�5�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �???????�?�?]t�E�?F]t�E�?��y��y�?�a�a�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���/hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@D         >                    �?Ly�'^��?Z           ��@               #                    �?~n��e�?z            @g@                                  �L@p�"�0�?a            �b@                                  �?�&=�w��?E            �Z@               
                   �b@�S����?
             3@                                  �J@�����H�?	             2@       ������������������������       �                     *@               	       
             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                   �K@���E�?;            �U@       ������������������������       �        8             U@                                  @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                      
             �?��V#�?            �E@                                 �r@X�<ݚ�?             2@                                   Q@      �?             (@                                  �?ףp=
�?	             $@                                  �M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                  pc@r�q��?             @                                  0v@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               "                    �?�J�4�?             9@                !       	          ����?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@        $       +                    @I@��+��?            �B@        %       &       
             �?"pc�
�?             &@        ������������������������       �                     �?        '       (                    Z@z�G�z�?             $@        ������������������������       �                     �?        )       *                    �B@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ,       =                   `c@$��m��?             :@       -       8                    �?�GN�z�?             6@       .       3                    �J@r�q��?             2@        /       2                    �?�q�q�?             @       0       1                    �I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        4       5                    �?�8��8��?	             (@       ������������������������       �                      @        6       7                   @_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        9       <       	             �?      �?             @       :       ;                   �\@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ?       �       
             �?�e&���?�           ��@       @       �                   �`@�K>��[�?$           �{@       A       �                    @M@6�I#r�?�             o@       B       k                    �?Te�$��?o             e@        C       L                   �f@�n_Y�K�?2            �S@        D       K                    �?\-��p�?             =@        E       J                   @_@      �?	             0@        F       G                    \@�q�q�?             @        ������������������������       �                     �?        H       I                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        
             *@        M       j                    �?Rg��J��?            �H@       N       _       	          ����?8�A�0��?             F@        O       P                    ]@p�ݯ��?             3@        ������������������������       �                     @        Q       V                   �^@     ��?
             0@        R       U                   �]@և���X�?             @       S       T                    �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        W       ^                   �e@�q�q�?             "@       X       ]       	          ����?؇���X�?             @       Y       \                    �?      �?             @       Z       [       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        `       i                   �q@�+e�X�?             9@       a       h       	             @ҳ�wY;�?             1@       b       c                   �\@������?
             .@        ������������������������       �                      @        d       e       	          ����?8�Z$���?             *@        ������������������������       �                      @        f       g                   j@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        l       o                   �Z@8�Z$���?=            �V@        m       n                   `_@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        p       q                   �h@������?7            �T@        ������������������������       �                     @@        r                           @L@�J�4�?#             I@       s       |       	             @�����H�?            �F@       t       y                    �?@4և���?             E@       u       v                    �?������?             B@       ������������������������       �                     A@        w       x                     H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        z       {                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        }       ~       	          ���@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	             �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �a@���(\��?3             T@       �       �                   �]@�n���?,             R@       �       �                   Pg@����?�?            �F@       ������������������������       �                     :@        �       �                    Y@�}�+r��?             3@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?PN��T'�?             ;@        �       �                    �?�q�q�?             (@       ������������������������       �                     @        �       �                   `@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                    �P@      �?              @       �       �                   �^@�q�q�?             @        ������������������������       �                      @        �       �       	          ����?      �?             @        ������������������������       �                     �?        �       �                   �d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @��(!i�?�            �h@       �       �                    �?X��t��?|             g@       �       �       	          ����?�.�?�P�?P             ^@        �       �                    @N@p�ݯ��?             3@       �       �                    @M@��S���?	             .@       �       �                    �?�n_Y�K�?             *@       �       �                   �n@      �?             $@       �       �                    X@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��'cy�?D            @Y@       �       �                   �b@�7��?5            �S@       �       �                   `a@@�E�x�?!            �H@        ������������������������       �                     .@        �       �                   �a@г�wY;�?             A@       �       �                   �b@P���Q�?             4@       ������������������������       �                     1@        �       �       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �f@ܷ��?��?             =@        �       �                   `U@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@        ������������������������       �                     7@        �       �                    �R@      �?,             P@       �       �                    �? ������?+            �O@       ������������������������       �        $            �J@        �       �                    n@ףp=
�?             $@       ������������������������       �                     @        �       �                   �n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?      �?             (@        ������������������������       �                     @        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �L@������?�            �q@       �       �                    �?:䠍[O�?�            @k@        �       �       	            �? 9�����?6             V@       �       �                   �b@�'N��?'            �N@       �       �       	             � 	��p�?             =@        ������������������������       �                      @        ������������������������       �                     ;@        �       �                   0f@     ��?             @@       �       �                   ``@
j*D>�?             :@       �       �                    �?      �?             4@        ������������������������       �                      @        �       �                    @G@�q�q�?             (@        �       �                   �c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   0m@�����H�?             ;@       ������������������������       �        
             1@        �       �                    @F@�z�G��?             $@        ������������������������       �                      @        �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �g@ ��WV�?[            @`@       �       �                    @L@0Ƭ!sĮ?Z             `@       �       �       	             @�Ń��̧?X            �_@       �       �                   @n@`o��b�?W             _@       ������������������������       �        5            �S@        �       �                    �?��<b�ƥ?"             G@       ������������������������       �                     =@        �       �                   @c@�IєX�?             1@        �       �                   �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                      @        �       �                   Hp@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �                         �a@��z4���?+            @Q@       �                          `P@�D����?             E@       �       �                    �?�������?             A@        �       �                   @`@      �?              @        ������������������������       �                     @        �       �                    �?z�G�z�?             @        �       �                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �                          �]@���B���?             :@        �       �       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                �_@�C��2(�?             6@                                 @N@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             ,@        ������������������������       �                      @                                 �?�<ݚ�?             ;@       ������������������������       �        	             0@        	                         a@�eP*L��?             &@       
            	          ����?����X�?             @        ������������������������       �                     �?                    	             �?r�q��?             @                                n@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B  ȫ�rV��?���T8�?��&�h��?v�e�]v�?�PM�\"�?�y���?tHM0���?�x+�R�?(������?^Cy�5�?�q�q�?�q�q�?      �?        333333�?�������?              �?      �?                      �?m��֡�?Ȥx�L��?      �?        UUUUUU�?UUUUUU�?              �?      �?        eMYS֔�?6eMYS��?�q�q�?r�q��?      �?      �?�������?�������?�������?�������?      �?                      �?              �?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?        �z�G��?{�G�z�?UUUUUU�?UUUUUU�?              �?      �?              �?        *�Y7�"�?�S�n�?/�袋.�?F]t�E�?      �?        �������?�������?              �?�q�q�?�q�q�?              �?      �?        vb'vb'�?�N��N��?]t�E�?�袋.��?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �(5�0�?�k�g��?K�p�ɵ�?��ㄍ��?a2�>�?h3�?R0�?8�Z$���?d���+��?ى�؉��?;�;��?�{a���?a����?      �?      �?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?                      �?              �??4և���?��S�r
�?颋.���?/�袋.�?Cy�5��?^Cy�5�?              �?      �?      �?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?              �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?      �?      �?      �?              �?      �?                      �?              �?      �?        R���Q�?���Q��?�������?�������?wwwwww�?�?              �?;�;��?;�;��?      �?        333333�?�������?              �?      �?                      �?      �?                      �?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?        ������?�|����?              �?{�G�z�?�z�G��?�q�q�?�q�q�?�$I�$I�?n۶m۶�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?      �?                      �?�����̼?ffffff�?r�qǱ?r�q��?l�l��?��I��I�?              �?(�����?�5��P�?�$I�$I�?۶m۶m�?              �?      �?                      �?h/�����?&���^B�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?4և��и?9/����?!Y�B�?����7��?wwwwww�?�?Cy�5��?^Cy�5�?�������?�?ى�؉��?;�;��?      �?      �?�������?UUUUUU�?              �?      �?                      �?              �?      �?                      �?��be�F�?`ҩy���?�A�A�?��[��[�?9/���?և���X�?              �?�?�?�������?ffffff�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?a���{�?��=���?      �?      �?              �?      �?                      �?              �?      �?      �?AA�?��}��}�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?              �?      �?              �?      �?        �v%jW��?��+Q��?��%�i?�?&�i?Y�?]t�E�?�E]t��?�����?ާ�d��?������?�{a���?              �?      �?              �?      �?;�;��?b'vb'v�?      �?      �?              �?�������?�������?�������?UUUUUU�?              �?      �?                      �?      �?              �?        �q�q�?�q�q�?              �?333333�?ffffff�?      �?              �?      �?      �?                      �?O��N���?;�;��?����?����?��<��<�?�a�a�?���{��?�B!��?      �?        ��7��M�?d!Y�B�?      �?        �?�?      �?      �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?̵s���?%~F���?�0�0�?z��y���?�������?�������?      �?      �?              �?�������?�������?      �?      �?              �?      �?              �?        ��؉���?ى�؉��?      �?      �?      �?                      �?]t�E�?F]t�E�?      �?      �?              �?      �?              �?                      �?�q�q�?9��8���?              �?t�E]t�?]t�E�?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��:hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�=         z                    �?�~8�e�?K           ��@              I       
             �?�n`���?C            @              >                   pt@��z��b�?�            �v@              ;                   �e@Pq�����?�            @u@              0                    @M@3u�cƵ?�            u@                                  Z@�f����?|             g@                                  @Y@���Q��?	             $@              	                    �?      �?              @        ������������������������       �                     �?        
                          0a@؇���X�?             @       ������������������������       �                     @                      
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @               /                   �a@XpBt,��?s            �e@                                 Pf@�'g�2�?\            �a@        ������������������������       �                     �J@                                    `@ףp=
�?<            �V@                                  �`@      �?             H@                                  �?      �?             8@        ������������������������       �                     @                                   �?@�0�!��?             1@                                  �?�θ�?
             *@                                   �I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �K@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        !       (       	          ����?؇���X�?             E@        "       #                    �H@X�<ݚ�?             "@        ������������������������       �                     @        $       '                    �?z�G�z�?             @       %       &                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        )       *                   @X@�FVQ&�?            �@@        ������������������������       �                     �?        +       .                    �?      �?             @@        ,       -                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                     @@        1       :       
             �?�"w����?_             c@        2       9                    �R@      �?             @@       3       8                    �O@�g�y��?             ?@       4       7                   @Z@@4և���?             ,@        5       6                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �        K             ^@        <       =                   @Z@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ?       H       	          ����?8����?             7@       @       E                    a@��
ц��?	             *@       A       D                   `]@����X�?             @        B       C                    ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        F       G                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        J       k       	          pff�?B��仱�?V            �`@       K       b                    �M@\`*�s�?:             U@       L       M                   `b@     ��?.             P@        ������������������������       �                     >@        N       U                   �c@�t����?             A@        O       P                    �?����X�?             @        ������������������������       �                     �?        Q       T                    �?r�q��?             @        R       S                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        V       a                    p@�+$�jP�?             ;@       W       X                    @C@�q�q�?             (@        ������������������������       �                      @        Y       Z                   @i@      �?	             $@        ������������������������       �                      @        [       \                    �D@      �?              @        ������������������������       �                     �?        ]       ^                     I@����X�?             @        ������������������������       �                     @        _       `                   @`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     .@        c       h                    V@��Q��?             4@        d       e                   �\@ףp=
�?             $@       ������������������������       �                      @        f       g                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        i       j                   �c@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        l       s                    �? \� ���?            �H@        m       n                   �V@D�n�3�?             3@        ������������������������       �                     @        o       r                    `@�8��8��?             (@        p       q                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        t       y                   `U@(;L]n�?             >@        u       v                    `@      �?              @       ������������������������       �                     @        w       x       	          033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             6@        {       �                    @L@ꀌ�N�?           `z@       |       �                    �?�2�MA��?�            �q@        }       �                   �p@      �?]             b@       ~                          `X@�eGk�T�?=            �W@        ������������������������       �                     �?        ������������������������       �        <            �W@        �       �       	          `ff�?ZՏ�m|�?             �H@       �       �                    �K@��Y��]�?            �D@       ������������������������       �                     C@        �       �       	          `ff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �r@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�f|��?]            �a@       �       �                   �Z@�8�So��?O            @^@        �       �       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   d@p/3�d��?L            �]@        �       �                    d@�eP*L��?             &@        �       �                    �G@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @z�G�z�?             @        ������������������������       �                     @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          `ff@�ʠ����?D            �Z@       �       �                   �z@0��_��?C            �Z@       �       �                    �?�#-���?B            @Z@        ������������������������       �                    �G@        �       �                   f@Riv����?+             M@       �       �                    �?�������?"             F@        ������������������������       �                     "@        �       �                   `p@��R[s�?            �A@       �       �       	          ����?ȵHPS!�?             :@       �       �       
             �?�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        �       �                   �f@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             ,@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @G@�GN�z�?             6@        ������������������������       �                     @        �       �                    �K@�X�<ݺ?             2@       ������������������������       �        	             ,@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @\@�����]�?N            �`@        �       �                    @N@ȵHPS!�?             :@        �       �                    �?      �?             @       �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `V@���7�?             6@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             4@        �       �       
             �?�A�|O��??            @[@       �       �                    �?4�	~���?'            @Q@       �       �       
             �?�K��&�?            �E@        �       �                    @؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �[@�q�q�?             B@        ������������������������       �                     @        �       �                    �?���!pc�?            �@@       �       �                    �?�ՙ/�?             5@       �       �                    ^@z�G�z�?	             .@        ������������������������       �                     �?        �       �                   c@؇���X�?             ,@        ������������������������       �                     @        �       �                   �c@      �?              @        ������������������������       �                     �?        �       �                   �c@؇���X�?             @        ������������������������       �                     @        �       �                   `\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    @�8��8��?             (@       �       �       	          ����?ףp=
�?             $@       �       �                   p`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @O@8�Z$���?             :@        ������������������������       �                     ,@        �       �                   �`@�q�q�?             (@        ������������������������       �                      @        �       �                   0`@z�G�z�?             $@        ������������������������       �                     @        �       �                     Q@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?z�G�z�?             D@       �       �                    �?�r����?             >@       �       �                   Pc@�J�4�?             9@       ������������������������       �        	             *@        �       �                    �?�q�q�?             (@        ������������������������       �                     @        �       �       	          ����?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �������?222222�?�c�1��?�9�s��?
V2k8�??������?�?~~~~~~�?��P�ʦ?����^��?���;��?��X��?�������?333333�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �>���T�?L�w�Z�?�^���?$T�ik��?              �?�������?�������?      �?      �?      �?      �?              �?�������?ZZZZZZ�?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?                      �?              �?�$I�$I�?۶m۶m�?�q�q�?r�q��?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        |���?>����?      �?              �?      �?      �?      �?              �?      �?                      �?              �?(�����?Cy�5��?      �?      �?�B!��?��{���?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        8��Moz�?d!Y�B�?�;�;�?�؉�؉�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?UUUUUU�?      �?                      �?              �?d\��?���7G��?��<��<�?b�a��?      �?      �?      �?        �������?�������?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?      �?      �?                      �?              �?/�����?B{	�%��?�������?�������?      �?              �?      �?              �?      �?      �?              �?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?              �?        ffffff�?�������?�������?�������?              �?      �?      �?              �?      �?        333333�?�������?      �?                      �?և���X�?
^N��)�?l(�����?(������?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �?�������?      �?      �?              �?      �?      �?              �?      �?                      �?�0�Y���?�oL���?��B���?6�����?      �?      �?��=�ĩ�?�X�0Ҏ�?              �?      �?        �>4և��?9/����?8��18�?������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �P}����?�^���?���#���?��!pc�?UUUUUU�?UUUUUU�?              �?      �?        ����c�?~ylE�p�?]t�E�?t�E]t�?UUUUUU�?�������?      �?                      �?�������?�������?      �?              �?      �?              �?      �?        �@�Ե�?7��XQ�?"5�x+��?�V�9�&�?�A�A�?_�_�?      �?        >�����?	�=����?t�E]t�?/�袋.�?      �?        X|�W|��?PuPu�?��N��N�?�؉�؉�?�Mozӛ�?d!Y�B�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?]t�E�?�袋.��?      �?        �q�q�?��8��8�?              �?      �?      �?              �?      �?        �)F�?$�\y@�?�؉�؉�?��N��N�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?�.�袋�?      �?      �?              �?      �?                      �?Y���%�?N��ش�?F��Q�g�?];0���?���)k��?��)kʚ�?۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?        t�E]t�?F]t�E�?�a�a�?�<��<��?�������?�������?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?�������?�������?      �?                      �?              �?              �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?              �?      �?        ffffff�?ffffff�?�������?�?�z�G��?{�G�z�?      �?        UUUUUU�?UUUUUU�?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        ffffff�?333333�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��5hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         �                    �?�&���?=           ��@              A                    �?нK���?C           ��@                      
             �?և���X�?�             k@                                  �?�p�I�?K            �]@                                  @a@
;&����?             7@                                  �?������?             .@       ������������������������       �                     &@        ������������������������       �                     @        	              	          `ff�?      �?              @        
              	          pff�?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                  pr@8��8���?>             X@                                 `_@Pq�����?7            @U@        ������������������������       �                    �E@                                   `@�����?             E@        ������������������������       �                     �?                      	          033�?��p\�?            �D@                      	          ����?@�0�!��?             1@       ������������������������       �        	             ,@        ������������������������       �                     @        ������������������������       �                     8@                                   �?�eP*L��?             &@                     	          ����?X�<ݚ�?             "@                     	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @               (                   �a@~	~���?=            �X@                !                    �L@ȵHPS!�?             J@       ������������������������       �                     ?@        "       #                   @]@����X�?
             5@        ������������������������       �                     @        $       '                   �]@�q�q�?             2@        %       &                    �?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        )       <                    �M@(옄��?!             G@       *       1                   Pc@�n_Y�K�?            �C@        +       0                   �b@      �?              @       ,       /                    �?���Q��?             @       -       .       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        2       ;                    �?¦	^_�?             ?@       3       :                   �_@H%u��?             9@        4       9                   �f@      �?             @       5       6                    �?      �?             @        ������������������������       �                      @        7       8                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        ������������������������       �                     @        =       @                   �_@؇���X�?             @        >       ?                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        B       �       
             �?H+��t��?�            �s@       C       v                   �b@ДXࣿ?�             q@       D       u                    �?`����?�            �o@       E       h                    �K@��S�ۿ?t            `h@       F       _                   pp@W�!?�?<            �X@       G       R                   `\@�X�C�?%             L@        H       O       	             @X�Cc�?	             ,@       I       J                    �?z�G�z�?             $@        ������������������������       �                      @        K       L                   @[@      �?              @       ������������������������       �                     @        M       N                   �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        P       Q       	             @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        S       X                   `b@�����?             E@       T       W                    �?      �?             @@        U       V       	             @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     <@        Y       ^                   `c@�z�G��?             $@        Z       [                    `@      �?             @        ������������������������       �                     �?        \       ]                    �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        `       g       	          ����? qP��B�?            �E@        a       b                   �Z@      �?              @        ������������������������       �                     @        c       d                    @H@      �?             @        ������������������������       �                      @        e       f                    @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �A@        i       t       	          ����?      �?8             X@        j       k       	          ����?�����H�?             ;@        ������������������������       �                     @        l       m                    @N@R���Q�?             4@        ������������������������       �                     "@        n       o       	          hff�?���!pc�?             &@        ������������������������       �                     �?        p       s                   �`@z�G�z�?             $@        q       r                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        '            @Q@        ������������������������       �                     �L@        w       x       	          433�?      �?             4@        ������������������������       �                     @        y       z       
             �?�t����?	             1@        ������������������������       �                     �?        {       |                   �`@      �?             0@        ������������������������       �                     @        }       ~                    q@z�G�z�?             $@       ������������������������       �                     @               �                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   a@v�X��?             F@       �       �                    �N@�5��?             ;@       �       �                    �?b�2�tk�?             2@        ������������������������       �                      @        �       �                    n@     ��?
             0@        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �a@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   pf@�t����?             1@       �       �                    �?      �?             0@        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     �?        �       �                    �?����?�            x@       �       �                    @�>4և��?�            @s@       �       �       
             �?������?�             q@        �       �                   �d@t�C�#��?2            �S@       �       �                   `X@TV����?%            �M@        ������������������������       �                     @        �       �                    �?\�����?$            �K@        �       �                   �^@�t����?             1@        �       �                   @q@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �^@ףp=
�?             $@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �N@�s��:��?             C@       �       �                     H@�	j*D�?             :@        ������������������������       �                     @        �       �       
             �?��<b���?             7@        ������������������������       �                      @        �       �                    �?؇���X�?             5@        �       �                   �h@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?      �?             0@        �       �       	          433�?�q�q�?             @       �       �                   pn@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �       �       	          `ff�?      �?	             (@       �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?R���Q�?             4@        �       �       	          ����?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �                   Pc@࿾��@�?�            `h@        �       �       	            �?�X����?             6@       ������������������������       �                     .@        ������������������������       �                     @        �       �       	            �?����� �?v            �e@       �       �                    �? ���?h             b@        �       �                    �?@4և���?             ,@        �       �                   pd@؇���X�?             @       ������������������������       �                     @        �       �                    f@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        ]            ``@        �       �       	          pff�? �Cc}�?             <@        ������������������������       �                     @        ������������������������       �                     9@        �       �       
             �?�ʻ����?             A@       �       �                    �?��Q��?             4@        �       �                   `@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �r@�t����?             1@       �       �                    p@z�G�z�?
             .@       �       �                   �j@�q�q�?             "@       ������������������������       �                     @        �       �                   `b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �B@؇���X�?	             ,@        ������������������������       �                     �?        �       �                    a@$�q-�?             *@        �       �                   �_@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@����?0            @S@       �       �       
             �?��.��?%            �N@       �       �                     P@���5��?!            �L@       �       �                    �J@HP�s��?             I@        �       �                   �`@����X�?             ,@        ������������������������       �                      @        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                   Pb@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     B@        �       �                   �j@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �f@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B�  \�\��?R��Q���?��S��?S�:+��?۶m۶m�?�$I�$I�?���?:�:��?Y�B��?�Mozӛ�?wwwwww�?�?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?�������?�������?�?~~~~~~�?              �?�a�a�?=��<���?      �?        ��+Q��?�]�ڕ��?�������?ZZZZZZ�?              �?      �?                      �?t�E]t�?]t�E�?�q�q�?r�q��?�������?�������?              �?      �?                      �?      �?        �)x9/�?h�����?��N��N�?�؉�؉�?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        ���,d�?ӛ���7�?;�;��?ى�؉��?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?��Zk���?�RJ)���?)\���(�?���Q��?      �?      �?      �?      �?              �?      �?      �?      �?                      �?      �?              �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?:�g *�?�	�Z��?������?�������?��i��i�?�eY�eY�?�?�������?1ogH�۹?�v���?%I�$I��?�m۶m��?�m۶m��?%I�$I��?�������?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�a�a�?=��<���?      �?      �?      �?      �?              �?      �?                      �?333333�?ffffff�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�}A_З?��}A�?      �?      �?              �?      �?      �?              �?      �?      �?      �?                      �?              �?      �?      �?�q�q�?�q�q�?              �?333333�?333333�?              �?t�E]t�?F]t�E�?      �?        �������?�������?      �?      �?      �?                      �?              �?              �?              �?      �?      �?      �?        �?<<<<<<�?              �?      �?      �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?颋.���?�.�袋�?/�����?h/�����?�8��8��?9��8���?              �?      �?      �?�q�q�?�q�q�?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?              �?�?<<<<<<�?      �?      �?      �?                      �?      �?        @��(C�?���y��?�$I�$I�?�m۶m��?�*alT�?T{N���?��td�@�?��7a~�?E�pR���?u_[4�?      �?        ߰�k��?A��)A�?�������?�������?۶m۶m�?�$I�$I�?      �?                      �?�������?�������?      �?      �?      �?                      �?      �?        �k(���?��k(��?;�;��?vb'vb'�?      �?        ��Moz��?��,d!�?      �?        �$I�$I�?۶m۶m�?�������?333333�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?      �?      �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        333333�?333333�?      �?      �?              �?      �?              �?        �1�1�?����?�E]t��?]t�E]�?      �?                      �?����B�?���"��?x����?����?|?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        %I�$I��?۶m۶m�?              �?      �?        �������?<<<<<<�?ffffff�?�������?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?�������?UUUUUU�?      �?                      �?      �?        �S{��?
qV~B��?������?�����?��Gp�?�}��?{�G�z�?q=
ףp�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?      �?                      �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@F         �       
             �?V�2���?7           ��@              g                   P`@�fC���?8           `@               J                    `@*T1e���?�             o@              E                    �?Z���c��?q            �g@              :       	          pff�?$�7�L��?S            �a@              #                    @J@�q�q�?<            �Y@                                   `r@�F�j��?            �J@                                 �p@X�<ݚ�?            �F@       	              	          ����?Hث3���?            �C@        
                           �?������?
             .@        ������������������������       �                     �?                      	          ����?d}h���?	             ,@                                  �?      �?             (@        ������������������������       �                     @                                   ]@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                    B@�q�q�?             8@        ������������������������       �                     @                                  �Q@�S����?
             3@        ������������������������       �                     �?                                   @D@�����H�?	             2@                                  0j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  pf@      �?             0@                                   �E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     @        !       "                   ({@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        $       9       	          ����?؇���X�?            �H@       %       .       	          ����?      �?             H@       &       -                    @L@`Jj��?             ?@        '       ,                   @d@8�Z$���?             *@       (       )                    �?�8��8��?             (@       ������������������������       �                     "@        *       +                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             2@        /       8                   @_@������?             1@       0       1                    �?     ��?
             0@        ������������������������       �                     �?        2       7                   �[@�r����?	             .@        3       4                   `_@�q�q�?             @        ������������������������       �                     @        5       6                     L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ;       >                   �\@$�q-�?            �C@        <       =       	          ���@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ?       @                   Pb@(;L]n�?             >@       ������������������������       �                     8@        A       B                    �?r�q��?             @        ������������������������       �                     @        C       D                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        F       G                    �? �q�q�?             H@       ������������������������       �                    �D@        H       I                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        K       \                    a@�0u��A�?&             N@       L       [                   �^@�S����?             C@       M       R                    �?V�a�� �?             =@        N       O       	          ����?z�G�z�?             @        ������������������������       �                     @        P       Q                   `[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       T                    @L@�8��8��?             8@        ������������������������       �                     $@        U       V                   �X@؇���X�?             ,@        ������������������������       �                     �?        W       Z                    �?$�q-�?             *@        X       Y                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     "@        ]       f                   �q@�GN�z�?             6@       ^       _       	          ����?��s����?             5@        ������������������������       �                      @        `       e                    @O@�KM�]�?             3@       a       b                    �?�X�<ݺ?
             2@       ������������������������       �                     0@        c       d                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        h       {                    �?`0�Ƒg�?�            �o@        i       p                    �?�T`�[k�?%            �J@       j       k                   �b@@-�_ .�?            �B@       ������������������������       �                     >@        l       m                   `a@����X�?             @        ������������������������       �                     �?        n       o                   xu@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        q       t                   pk@      �?
             0@        r       s                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        u       z                   �e@"pc�
�?             &@       v       y                   �b@ףp=
�?             $@        w       x       	          ����?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        |       �                    @��(\���?|             i@       }       �                   �u@ �r�ɻ?w            �g@       ~       �                   �b@p��D��?s             g@              �                    �?�|1)�?@            �Z@        �       �       	          033�?r�q��?             (@       �       �                    �H@�C��2(�?             &@        �       �                     H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   h@��K2��?9            �W@        �       �                     M@h�����?             <@        �       �                   @a@�C��2(�?             &@       ������������������������       �                     "@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             1@        ������������������������       �        )            �P@        �       �                   �b@l{��b��?3            �S@        �       �                    �N@\-��p�?             =@       �       �                   �_@      �?             0@       ������������������������       �                      @        �       �                   �a@      �?              @       �       �                    �?z�G�z�?             @       �       �                    `@�q�q�?             @        ������������������������       �                     �?        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        �       �                    �Q@`2U0*��?             I@       �       �                    �?@��8��?             H@       ������������������������       �                    �D@        �       �       	             �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                     O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    b@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@0��k���?�             z@       �       �                   @E@�3��r�?�            `q@        �       �                    �?�d�����?             3@       �       �                   `\@@4և���?	             ,@        �       �                   �X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?8L�0�h�?�            0p@        �       �       	          pff�?�GN�z�?             F@       �       �                    �?(N:!���?            �A@       �       �                    �?H%u��?             9@       �       �                    �?��2(&�?             6@        ������������������������       �                     $@        �       �                    �D@      �?	             (@        ������������������������       �                     @        �       �                   �p@�q�q�?             "@        ������������������������       �                     @        �       �                   �r@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                     C@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �n@�q�q�?             "@       �       �                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �? �LV�-�?�            �j@       �       �                    �?@��d�`�?             i@        �       �       	          433�? 7���B�?             ;@       ������������������������       �                     7@        �       �                   0a@      �?             @        �       �                   pg@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        i            �e@        �       �       	          033�?�r����?	             .@       �       �                    �?@4և���?             ,@        �       �                    �I@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        �                          �?��c:�?N            @a@       �       �                    �?�B�����?;             Z@        �       �                   @V@     ��?             @@        ������������������������       �                     @        �       �                   �d@ 	��p�?             =@       ������������������������       �                     4@        �       �                   0r@�<ݚ�?             "@       ������������������������       �                     @        �       �                   @_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �N@*O���?)             R@       �       �                    �M@�G��l��?             E@       �       �                   @]@�P�*�?             ?@        ������������������������       �                     @        �       �                    a@r�q��?             8@        �       �       	          ����?8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �L@"pc�
�?             &@        �       �       	          ����?���Q��?             @       �       �                    c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   P`@���|���?             &@        ������������������������       �                     @        �       �       	          @33�?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @                     	          `ff�?z�G�z�?             >@                                �?�nkK�?             7@        ������������������������       �                     *@                                  P@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@                                `c@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        	      
                   �?������?             A@        ������������������������       �                      @                                 �?     ��?             @@                                S@��+7��?             7@                    	             �?և���X�?             @                                [@���Q��?             @        ������������������������       �                      @                                �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                �q@      �?	             0@       ������������������������       �                     "@                                  O@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  � ���Y�?�o�6S�?VD�Tw��?�.�*�S�?p���?�#�9�?��i��i�?Y�eY�e�?C��X��?^���S��?UUUUUU�?UUUUUU�?��sHM�?:�&oe�?�q�q�?r�q��?�i�i�?��-��-�?�?wwwwww�?      �?        ۶m۶m�?I�$I�$�?      �?      �?              �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?(������?^Cy�5�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?�B!��?���{��?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�?xxxxxx�?      �?      �?      �?        �?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?        ;�;��?�؉�؉�?�q�q�?9��8���?              �?      �?        �?�������?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?UUUUUU�?�������?              �?�$I�$I�?�m۶m��?      �?                      �?�������?�������?^Cy�5�?(������?a���{�?��{a�?�������?�������?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�袋.��?]t�E�?z��y���?�a�a�?              �?�k(���?(�����?��8��8�?�q�q�?      �?              �?      �?              �?      �?                      �?              �?����Q�?&b�C���?"5�x+��?���!5��?к����?S�n0E�?              �?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?              �?      �?�������?�������?      �?                      �?/�袋.�?F]t�E�?�������?�������?      �?      �?      �?                      �?      �?                      �?333333�?�������?o��2�|�?�ќ5(�?����y�?�cxq�?"5�x+��?W�9�&�?UUUUUU�?�������?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        W�+�Ʌ?��Q�٨�?�$I�$I�?�m۶m��?F]t�E�?]t�E�?              �?      �?      �?              �?      �?                      �?              �?�&��jq�?${�ґ�?�{a���?a����?      �?      �?              �?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?              �?{�G�z�?���Q��?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?r�q��?              �?      �?        �؉�؉�?��؉���?W��_��?Le{�ݸ?y�5���?Cy�5��?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?�������?�������?      �?                      �?M�]��d�?.�!J粩?�袋.��?]t�E�?|�W|�W�?�A�A�?)\���(�?���Q��?��.���?t�E]t�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?      �?              �?        �������?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?��i���?X:Ɂ���?ףp=
��?{�G�zt?	�%����?h/�����?      �?              �?      �?      �?      �?      �?                      �?      �?              �?        �������?�?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?-d!Y��?�7��Mo�?b'vb'v�?;�;��?      �?      �?              �?������?�{a���?      �?        9��8���?�q�q�?      �?              �?      �?      �?                      �?�q�q�?�q�q�?1�0��?��y��y�?�RJ)���?�Zk����?      �?        UUUUUU�?UUUUUU�?;�;��?;�;��?      �?                      �?/�袋.�?F]t�E�?333333�?�������?      �?      �?      �?                      �?      �?              �?        F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?              �?      �?        �������?�������?�Mozӛ�?d!Y�B�?      �?        �������?�������?              �?      �?        �$I�$I�?�m۶m��?              �?      �?        �?xxxxxx�?      �?              �?      �?Y�B��?zӛ����?�$I�$I�?۶m۶m�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?�$I�$I�?�m۶m��?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJJ�/xhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�C         �                   �b@�lb���?;           ��@              }       
             �?m��1��?�           ��@              V                   P`@\�1���?           �z@                                   �?�����?�            �l@                                   �?b�2�tk�?             B@                                 h@ҳ�wY;�?             A@        ������������������������       �                     @                                   @I@և���X�?             <@        	       
                    Z@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@                                   �?b�2�tk�?             2@        ������������������������       �                     @                                  (s@d}h���?	             ,@                                 �^@8�Z$���?             *@                                  @q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  hq@�C��2(�?             &@        ������������������������       �                     @                                   �?z�G�z�?             @                                  �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                  �U@ی�
��?o            @h@        ������������������������       �                      @               =                   �^@�8��8��?n             h@              ,                    �?���Ls�?I            @`@                '                    �O@�X����?             6@       !       "       
             �?ףp=
�?             $@        ������������������������       �                      @        #       &                   �l@      �?              @        $       %                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        (       )                   `X@      �?             (@        ������������������������       �                     @        *       +                    �P@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        -       2       	          @33�?X'"7��?:             [@        .       1                   `X@l��\��?             A@        /       0                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ;@        3       <                   �[@�?�|�?&            �R@        4       5                   �Z@ >�֕�?            �A@        ������������������������       �                     0@        6       7                   ph@�KM�]�?             3@        ������������������������       �                      @        8       9                   Pk@"pc�
�?             &@        ������������������������       �                     �?        :       ;       	             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                    �C@        >       A       
             �?t�7��?%             O@        ?       @                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        B       Q                    `@���5��?"            �L@        C       P                    �?����X�?             5@       D       K                    �?      �?             0@        E       F                    �?؇���X�?             @        ������������������������       �                     �?        G       H                   @k@r�q��?             @        ������������������������       �                     @        I       J                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        L       M                   8p@X�<ݚ�?             "@        ������������������������       �                     @        N       O                   �p@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        R       S                    �?������?             B@       ������������������������       �                     >@        T       U                     N@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        W       x                    @�����?�            �h@       X       q                   @s@ �r�ѷ?|             g@       Y       l                   `f@�{���l�?n            �c@       Z       [                   �j@�'F�3�?j            �b@       ������������������������       �        6            �S@        \       ]                    k@0z�(>��?4            �Q@        ������������������������       �                     �?        ^       k                   Pa@��?^�k�?3            �Q@       _       j                    �?�nkK�?#             G@       `       i       	          ����? 	��p�?             =@        a       f                    �?8�Z$���?             *@       b       e                    b@�C��2(�?	             &@        c       d                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        g       h       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     1@        ������������������������       �                     8@        m       p                   �a@      �?              @        n       o                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        r       w                    �Q@�+$�jP�?             ;@       s       v                    �?H%u��?             9@        t       u                    w@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             0@        ������������������������       �                      @        y       z                   l@�	j*D�?             *@        ������������������������       �                      @        {       |                    �L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                    �?je�24�?~            �h@              �                   @E@H�ՠ&��?d            @d@        �       �       	            �?��
ц��?             :@       �       �                    @D@z�G�z�?	             .@        ������������������������       �                     �?        �       �                    �?؇���X�?             ,@       �       �                    ^@$�q-�?             *@       ������������������������       �                     $@        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?�wY;��?U             a@        �       �                   �b@      �?             4@       �       �                   �e@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �        
             *@        �       �                   p`@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       	             �? _�@�Y�?H             ]@       �       �       	            �?�H�I���?F            @\@       ������������������������       �        =            @Y@        �       �                   0p@�8��8��?	             (@       ������������������������       �                     $@        �       �                   pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   Pa@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?^������?            �A@       �       �       	          hff�?      �?             8@        �       �                    �?�<ݚ�?             "@       �       �                   e@����X�?             @       �       �                     P@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�q�q�?
             .@       �       �                    S@r�q��?             (@        �       �       	             �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �       �                    �?>���?�            `r@        �       �                    �?�O�w���?;            �V@       �       �                   �r@�O�y���?0            �R@       �       �                   pn@�0u��A�?(             N@       �       �                   @^@�ʻ����?             A@        �       �                   d@      �?              @       ������������������������       �                     @        �       �                   pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   l@�	j*D�?             :@       �       �                   `a@���Q��?
             4@       �       �       
             �?z�G�z�?             .@        ������������������������       �                     �?        �       �                   �_@؇���X�?             ,@        �       �                    _@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?8�Z$���?             :@        �       �                   pc@$�q-�?	             *@        �       �       	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          @33�?�θ�?	             *@       �       �                    �?և���X�?             @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?������?             .@       �       �                   �d@ףp=
�?             $@       ������������������������       �                     @        �       �                   0e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     0@        �       �       
             �?|g�&��?{            `i@        �       �                    �?Np�����?             �I@        �       �                    �?      �?
             0@       ������������������������       �                     $@        �       �                   �b@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �f@">�֕�?            �A@       �       �                     F@      �?             @@        �       �                   �l@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �L@8�Z$���?             :@        �       �                    �?�z�G��?             $@        ������������������������       �                      @        �       �                   e@      �?              @       ������������������������       �                     @        �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             0@       �       �                     O@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �_@p�|�i�?[             c@        �       �                   pn@0�z��?�?#             O@        �       �                    @G@���7�?             6@       ������������������������       �                     1@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     D@        �                         `@�X�<ݺ?8            �V@                                  �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @              
                   @ 7���B�?5            @T@             	                  �c@�?�|�?/            �R@                                `a@8�Z$���?	             *@        ������������������������       �                     @                                �c@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        &            �N@                                �k@؇���X�?             @                    	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  �y�@$�?�4æ�m�?��؉���?;�;��?|�g��?� [8��?���(�?�T>��u�?�8��8��?9��8���?�������?�������?      �?        �$I�$I�?۶m۶m�?�������?�������?              �?      �?        9��8���?�8��8��?      �?        ۶m۶m�?I�$I�$�?;�;��?;�;��?      �?      �?      �?                      �?F]t�E�?]t�E�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�Q�/�~�?��tT��?      �?        �������?�����*�?z�z��?�����?]t�E]�?�E]t��?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?B{	�%��?Lh/����?�������?------�?۶m۶m�?�$I�$I�?              �?      �?                      �?к����?*�Y7�"�?�A�A�?��+��+�?              �?(�����?�k(���?              �?F]t�E�?/�袋.�?      �?        �������?�������?      �?                      �?              �?��Zk���?SJ)��R�?�������?�������?      �?                      �?��Gp�?�}��?�$I�$I�?�m۶m��?      �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        r�q��?�q�q�?              �?�������?UUUUUU�?      �?                      �?              �?�q�q�?�q�q�?              �?UUUUUU�?�������?              �?      �?        �����?/,FBi��?��,d!�?�7��Mo�?Kz���?�-4`I/�?��c.��?��v[�?              �?H���@��?�ԓ�ۥ�?      �?        �A�A�?_�_��?d!Y�B�?�Mozӛ�?�{a���?������?;�;��?;�;��?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?                      �?              �?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?B{	�%��?/�����?���Q��?)\���(�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ;�;��?vb'vb'�?              �?�������?�������?              �?      �?        ���P��?8�ӹ���?������?{	�%���?�؉�؉�?�;�;�?�������?�������?              �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?ZZZZZZ�?ZZZZZZ�?      �?      �?n۶m۶�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        #,�4�r�?�{a���?x�!���?x�!���?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?_�_��?uPuP�?      �?      �?9��8���?�q�q�?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?�������?333333�?              �?      �?                      �?      �?                      �?��+�P�?��E�_�?�~�~��?�@�@�?�6�i�?~��K~�?�������?�������?�������?<<<<<<�?      �?      �?              �?      �?      �?      �?                      �?vb'vb'�?;�;��?333333�?�������?�������?�������?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ;�;��?;�;��?;�;��?�؉�؉�?�������?�������?              �?      �?                      �?�؉�؉�?ى�؉��?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?wwwwww�?�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?              �?      �?                      �?��v���?��%f-�?______�?PPPPPP�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�A�A�?_�_��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?333333�?ffffff�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?      �?        �k(����?^Cy�5�?|���{�?�B!��?�.�袋�?F]t�E�?      �?        �������?�������?      �?                      �?      �?        ��8��8�?�q�q�?9��8���?�q�q�?      �?                      �?	�%����?h/�����?*�Y7�"�?к����?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���WhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@>         �       
             �?:���sQ�?:           ��@              E                    �?�paRC4�?M            �@                                  �?�-���i�?�            pw@                                   �N@`��}3��?            �J@                                  �L@�'�=z��?            �@@                     	          ����?�n_Y�K�?             :@                                 @c@�	j*D�?	             *@              	                    @I@      �?             (@       ������������������������       �                     @        
                           �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                  ``@$�q-�?             *@                                  h@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@                                  Pa@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                      	          ����?P���Q�?
             4@                                  @O@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     $@                                  �U@�nkK�?�             t@        ������������������������       �                     �?               "                    Z@����<�?�            t@                                  �a@�<ݚ�?             "@       ������������������������       �                     @                !                    �I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        #       $                    �?@o-4j�?�            �s@        ������������������������       �        !             M@        %       0                    �?`n�:�6�?�            �o@        &       '       	          ����?�8��8��?+             N@       ������������������������       �                     A@        (       /                    �M@���B���?             :@       )       .       	          ����?�eP*L��?	             &@       *       -                    b@r�q��?             @       +       ,                    a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@        1       2                   Pe@��4+̰�?t            @h@        ������������������������       �        #            �P@        3       B                   0c@     �?Q             `@       4       5                   �e@`�c�г?N             _@        ������������������������       �                      @        6       A                   �a@ ;=֦��?M            �^@       7       @                   �\@p�|�i�?/             S@        8       9       	             �?�θ�?
             *@        ������������������������       �                     �?        :       ;                   �j@r�q��?	             (@        ������������������������       �                     �?        <       =                    @J@�C��2(�?             &@        ������������������������       �                     @        >       ?                     K@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        %            �O@        ������������������������       �                     G@        C       D                   `c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        F       o                   `_@��l�\��?g             e@        G       V                   �a@=��T�?-            �Q@        H       S                    @P@8����?             7@       I       R       	             �?r�q��?             2@        J       Q                   �_@      �?              @       K       P                    �?r�q��?             @       L       M                    @K@      �?             @        ������������������������       �                      @        N       O                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        T       U                   `]@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        W       X                   @J@��|�5��?            �G@        ������������������������       �                     @        Y       Z                   �Q@"pc�
�?             F@        ������������������������       �                      @        [       n                    �?؇���X�?             E@       \       e                    �?ףp=
�?             D@        ]       ^                   Pl@      �?             (@        ������������������������       �                     @        _       `                    �I@���Q��?             @        ������������������������       �                      @        a       b       	             �?�q�q�?             @        ������������������������       �                     �?        c       d                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       m                    �H@h�����?             <@        g       l                    ]@@4և���?             ,@        h       k                   pf@r�q��?             @       i       j       	          @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        	             ,@        ������������������������       �                      @        p       w                    @H@J����?:            �X@        q       r                    �?�����?	             3@        ������������������������       �                     @        s       t       	          433�?��
ц��?             *@        ������������������������       �                     @        u       v                    �E@      �?              @        ������������������������       �                      @        ������������������������       �                     @        x       �                    f@�Q��k�?1             T@       y       �                   �e@��|��?0            �S@       z                           �?��(�2Y�?-            �R@        {       ~       	          `ff�?���Q��?             $@       |       }                   �o@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?     �?&             P@        �       �                     L@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @N@XB���?#             M@       ������������������������       �                     C@        �       �       	          `ff�?ףp=
�?             4@       �       �                    @z�G�z�?             $@       �       �                    b@�����H�?             "@        ������������������������       �                     @        �       �                    �O@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �       	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @E@p�~;��?�            `w@        �       �                    �?�%^�?            �E@       �       �                    �?8^s]e�?             =@        �       �       	          -33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?l��
I��?             ;@        �       �                     F@�q�q�?             (@        ������������������������       �                     �?        �       �       	          433�?���!pc�?             &@        ������������������������       �                     @        �       �                   `@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             .@        �       �                    �?؇���X�?             ,@       �       �                     F@�8��8��?             (@        �       �                    @D@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�j1;#j�?�            �t@        �       �                    �?<=�,S��?,            �Q@       �       �                    @L@������?!            �I@       �       �                    �? �Cc}�?             <@        �       �                   �^@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        �       �                   0k@�û��|�?             7@        ������������������������       �                     @        �       �                   �c@�\��N��?             3@        ������������������������       �                     @        �       �                    @�	j*D�?             *@       �       �                    �L@"pc�
�?             &@        �       �                   0d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �N@�����H�?             "@       ������������������������       �                     @        �       �                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    n@�d�����?             3@        �       �       	          ����?      �?             @        ������������������������       �                      @        �       �                   `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�r����?             .@        ������������������������       �                      @        ������������������������       �                     *@        �       �       	          pff�?���(`�?�            Pp@       �       �                   �c@�߄��i�?�            �l@       �       �                    @L@ aqk+�?T            `a@       �       �                    �?�6H�Z�?D            @]@       ������������������������       �        2            �U@        �       �                   `b@(;L]n�?             >@       ������������������������       �                     9@        �       �                   c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    _@���7�?             6@        �       �                    @M@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                   Pd@ףp=
�?:            �V@        �       �                    �?����X�?             <@        ������������������������       �                     @        �       �                    a@���N8�?             5@       ������������������������       �        	             .@        �       �                    �?r�q��?             @       �       �                    d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �f@0�z��?�?)             O@       ������������������������       �        "            �I@        �       �                   @b@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                    �?     ��?             @@        ������������������������       �                     @        �       �                   �_@      �?             :@        ������������������������       �                     @        �       �                    �?8�A�0��?             6@       �       �                     M@      �?             0@       ������������������������       �                     "@        �       �                    �?և���X�?             @       �       �                    @�q�q�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �p@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  q���7T�?Ȏ �U�?�������?�?�{ͅ�)�?�PFo�Z�?M0��>��?�琚`��?|���?|��|�?ى�؉��?;�;��?vb'vb'�?;�;��?      �?      �?      �?        �������?333333�?              �?      �?                      �?;�;��?�؉�؉�?      �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?                      �?�������?ffffff�?�������?�������?      �?                      �?              �?d!Y�B�?�Mozӛ�?      �?        ��;6��?3�O�<��?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?� � �?�-��-��?              �?��b�X,�?���t:��?UUUUUU�?UUUUUU�?              �?ى�؉��?��؉���?]t�E�?t�E]t�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �? tT����?_\����?              �?      �?     ��?��RJ)��?��Zk���?      �?        XG��).�?�%C��6�?^Cy�5�?�k(����?�؉�؉�?ى�؉��?      �?        UUUUUU�?�������?      �?        F]t�E�?]t�E�?              �?UUUUUU�?�������?      �?                      �?              �?              �?      �?      �?      �?                      �?ƵHPS!�?��WV��?�:��:��?�������?8��Moz�?d!Y�B�?UUUUUU�?�������?      �?      �?UUUUUU�?�������?      �?      �?              �?      �?      �?      �?                      �?              �?      �?                      �?�������?�������?      �?                      �?br1���?x6�;��?              �?/�袋.�?F]t�E�?              �?۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�m۶m��?�$I�$I�?n۶m۶�?�$I�$I�?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?                      �?z;Cb���?Cb�ΐ��?Q^Cy��?^Cy�5�?      �?        �;�;�?�؉�؉�?      �?              �?      �?      �?                      �?�������?�������?� � �?˷|˷|�?*�Y7�"�?�����?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?     ��?UUUUUU�?�������?      �?                      �?�{a���?GX�i���?              �?�������?�������?�������?�������?�q�q�?�q�q�?              �?�������?�������?      �?                      �?      �?                      �?      �?      �?              �?      �?              �?        �X͞���?�ʄm�?�}A_�?�}A_��?	�=����?|a���?      �?      �?      �?                      �?h/�����?Lh/����?UUUUUU�?UUUUUU�?              �?F]t�E�?t�E]t�?      �?              �?      �?              �?      �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?      �?              �?      �?        '�쪉*�?eWMT�U�?�A�A�?X|�W|��?xxxxxx�?�?%I�$I��?۶m۶m�?      �?      �?              �?      �?              �?        8��Moz�?��,d!�?      �?        y�5���?�5��P�?      �?        ;�;��?vb'vb'�?F]t�E�?/�袋.�?      �?      �?      �?                      �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        y�5���?Cy�5��?      �?      �?      �?              �?      �?      �?                      �?�?�������?      �?                      �?g��o��?Ȥx�L��?&��pv�?��w���?O�&!��?4,�T�w�?�������?���?      �?        �������?�?      �?        �������?�������?              �?      �?        �.�袋�?F]t�E�?۶m۶m�?�$I�$I�?              �?      �?              �?        �������?�������?�m۶m��?�$I�$I�?              �?��y��y�?�a�a�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?        |���{�?�B!��?      �?        ]t�E�?F]t�E�?      �?                      �?      �?      �?      �?              �?      �?              �?颋.���?/�袋.�?      �?      �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?�������?              �?      �?        �t�bub�o=     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         �                    �?�s����?E           ��@              G                    �?NQ����?[           �@                                   �?.}Z*�?�            �j@               	                    �E@�99lMt�?            �C@                                  �V@z�G�z�?             @        ������������������������       �                     @                      
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        
                          pc@�t����?             A@                                 �`@8�A�0��?             6@                                  �?�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @                                   �M@�8��8��?             (@       ������������������������       �                     "@                                  �t@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               *       
             �?l�Ӑ���?p            �e@              %                   pr@@��j$޷?B            �Y@                     
             �?��V�I��?<            �W@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               $                    �?p�C��?9            �V@                      	          ����?���7�?             F@       ������������������������       �                     5@                      	          ����?���}<S�?             7@        ������������������������       �                     �?                !                   �k@���7�?             6@        ������������������������       �                     *@        "       #                   �k@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �G@        &       '                   �]@      �?              @        ������������������������       �                     @        (       )                    �G@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        +       @                    �?�q�q�?.             R@       ,       ;                   �_@�<ݚ�?'            �O@       -       :       	          833�?X�<ݚ�?             ;@       .       9                   �q@�LQ�1	�?             7@       /       4                   �b@���y4F�?             3@       0       1       	          ����?$�q-�?
             *@       ������������������������       �                     &@        2       3                    V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        5       8                   Pl@      �?             @       6       7                   �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        <       =                   �c@�X�<ݺ?             B@       ������������������������       �                     7@        >       ?                   �j@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        A       F                    @J@�<ݚ�?             "@       B       C       	          ,33ӿ�q�q�?             @        ������������������������       �                     @        D       E                   `\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        H       g                    �?�GT����?�            �t@        I       X       
             �?h���J;�?f            �c@        J       Q                   l@�q�����?             9@        K       P                    �K@z�G�z�?             $@       L       O                   @_@�q�q�?             @        M       N                    �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        R       W                   �`@�q�q�?
             .@       S       T                    �?r�q��?             (@        ������������������������       �                     @        U       V                    �I@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        Y       `                    �?�5[|/��?W            �`@        Z       [                   �p@���Q��?             .@       ������������������������       �                      @        \       _                   �f@؇���X�?             @       ]       ^                    d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        a       b                    @L@�6H�Z�?O            @]@       ������������������������       �        G            @Y@        c       d       	          ����?      �?             0@       ������������������������       �                     *@        e       f                    �M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        h       �       
             �?B0�8���?m            �e@        i       j                    @F@R_u^|�?-            �Q@        ������������������������       �                     &@        k       t       	          ����?�q�q�?'             N@        l       s                    �?�����?             5@        m       r                   �Z@�<ݚ�?             "@       n       o                    \@�q�q�?             @        ������������������������       �                      @        p       q                   0a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        u       v       	          833�?��
ц��?            �C@        ������������������������       �                      @        w       z                    �?��J�fj�?            �B@        x       y                   �Z@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        {       |       
             �?d��0u��?             >@        ������������������������       �                     @        }       �                    �?l��
I��?             ;@       ~                           �K@��S���?	             .@        ������������������������       �                     @        �       �                    �Q@�z�G��?             $@       �       �                   c@      �?              @        ������������������������       �                     @        �       �                    @�q�q�?             @        ������������������������       �                     �?        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �       	             @ȵHPS!�?@             Z@       �       �                    �?h�a��?=            @X@        �       �                    �Q@�8��8��?             B@       ������������������������       �                    �@@        ������������������������       �                     @        �       �                   `X@�]0��<�?'            �N@        ������������������������       �                     �?        �       �                    `@ �.�?Ƞ?&             N@        �       �                    _@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        "            �J@        ������������������������       �                     @        �       �                   �b@&�X~v��?�            Pw@       �       �                    �?������?�            pt@       �       �                    �L@     ��?�             p@       �       �                   �m@P��-�?[            �c@       �       �                    �?Df/��?7            �W@       �       �                    @K@z�G�z�?'            @P@       �       �       	             �?ZՏ�m|�?            �H@        ������������������������       �                     "@        �       �                   �m@z�G�z�?             D@       �       �                   �W@$G$n��?            �B@        ������������������������       �                     �?        �       �       	             �?�����H�?             B@       �       �                   0a@z�G�z�?             4@       �       �                    `@�t����?	             1@       �       �                   �a@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �h@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �i@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             0@        ������������������������       �                     @        �       �                   �d@     ��?             0@        ������������������������       �                      @        �       �                   �[@      �?              @        ������������������������       �                     @        �       �                   �`@      �?             @        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@        �       �                    �?�i�y�?$            �O@        �       �                   @_@�<ݚ�?             "@        �       �                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   0`@؇���X�?             @        �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     K@        �       �                   �Z@��F�D�?L            �X@        �       �                    �O@P���Q�?             4@       ������������������������       �        	             (@        �       �                     P@      �?              @        �       �                   �Y@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@�Fǌ��?<            �S@       ������������������������       �        ,            �K@        �       �                   �`@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        �       �                   b@�Y�R_�?&            �Q@       �       �       
             �?����"�?              M@       �       �                   �`@8����?             G@       �       �       	          033�?�t����?             A@       �       �                   �q@���y4F�?             3@       �       �                    �?�t����?             1@        ������������������������       �                     @        �       �                     P@8�Z$���?	             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             .@        �       �       	             �?r�q��?             (@        ������������������������       �                     �?        �       �                    �?�C��2(�?             &@       ������������������������       �                     @        �       �                   �a@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@        �       �       
             �?
;&����?             G@        �       �                   `a@�d�����?             3@       �       �                    @E@      �?             $@       �       �       	             �?r�q��?             @        �       �                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?��}*_��?             ;@        ������������������������       �                     "@        �       �                   @`@X�<ݚ�?             2@       �       �                   `Z@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �e@���|���?             &@       �       �       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��mQ��?-I׺��?KA����?k}U
���?�
��V�?�z2~���?5H�4H��?�o��o��?�������?�������?              �?      �?      �?              �?      �?        �������?�������?颋.���?/�袋.�?�������?�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        /�I���?�7[�~��?�?nnnnnn�?AL� &W�?<�����?UUUUUU�?UUUUUU�?      �?                      �?h�h��?��K��K�?F]t�E�?�.�袋�?              �?d!Y�B�?ӛ���7�?      �?        F]t�E�?�.�袋�?              �?�q�q�?�q�q�?      �?                      �?              �?      �?      �?              �?�������?333333�?              �?      �?        �������?�������?9��8���?�q�q�?r�q��?�q�q�?Nozӛ��?d!Y�B�?6��P^C�?(������?�؉�؉�?;�;��?      �?              �?      �?              �?      �?              �?      �?      �?      �?              �?      �?                      �?              �?              �?��8��8�?�q�q�?      �?        ;�;��?;�;��?              �?      �?        �q�q�?9��8���?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?l��(�?P�M�_�?����� �?9A���?�p=
ף�?���Q��?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        N6�d�M�?'�l��&�?333333�?�������?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?���?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �JC�}�?��jyc�?2~�ԓ��?�@�6�?      �?        UUUUUU�?UUUUUU�?�a�a�?=��<���?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?              �?�؉�؉�?�;�;�?      �?        к����?�"�u�)�?�m۶m��?�$I�$I�?              �?      �?        wwwwww�?DDDDDD�?      �?        h/�����?Lh/����?�?�������?      �?        333333�?ffffff�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?��N��N�?�؉�؉�?�D�a�Y�?���Id�?UUUUUU�?UUUUUU�?      �?                      �?\2�h��?;ڼOqɠ?              �?wwwwww�?�?۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?�?�����?0�J��?���]8��?��A��.�?      �?     ��?R��fu�?6��(S��?G}g����?� &W��?�������?�������?9/����?�>4և��?              �?�������?�������?���L�?к����?      �?        �q�q�?�q�q�?�������?�������?�?<<<<<<�?�q�q�?9��8���?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?              �?      �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?              �?AA�?�������?�q�q�?9��8���?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?[�R�֯�?j�J�Z�?�������?ffffff�?              �?      �?      �?      �?      �?              �?      �?                      �?�3���?1���M��?              �?UUUUUU�?�������?      �?                      �?�z2~���?���@��?�i��F�?	�=����?8��Moz�?d!Y�B�?�?<<<<<<�?(������?6��P^C�?�?<<<<<<�?              �?;�;��?;�;��?              �?      �?              �?                      �?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?        �������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�Mozӛ�?Y�B��?y�5���?Cy�5��?      �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?_B{	�%�?B{	�%��?      �?        �q�q�?r�q��?�$I�$I�?۶m۶m�?      �?                      �?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��khG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�C         �                    �?\r��ۖ�?E           ��@              S       
             �?^�L�8�?N           0�@               <                   ``@     8�?v             h@                                  @K@�D����?N            �_@                     	          ����?�p����?)            �N@                                   �? �o_��?             9@       ������������������������       �                     .@               	                    @E@�z�G��?             $@        ������������������������       �                     @        
                           �?      �?             @        ������������������������       �                     @        ������������������������       �                     @                                   �?      �?             B@                                   �?��
ц��?             *@        ������������������������       �                     @        ������������������������       �                     @                                  �[@���}<S�?             7@                                  Pi@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                      	          ���@���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?               /                    @O@��&����?%            @P@                     	          ���ٿ���H��?             E@        ������������������������       �                     @                      
             �?؇���X�?            �A@                                  �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               .                    �?<���D�?            �@@               #                   `X@PN��T'�?             ;@        !       "                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       -                    @H%u��?             9@       %       &                    �L@�8��8��?             8@        ������������������������       �                     ,@        '       ,                    l@z�G�z�?             $@       (       )       	          ����?�q�q�?             @        ������������������������       �                      @        *       +                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        0       ;                   �{@
;&����?             7@       1       8                   `@�G�z��?             4@        2       7                    �?�q�q�?             (@        3       6                   @_@z�G�z�?             @       4       5                   @d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        9       :                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        =       B       
             �?"pc�
�?(            �P@        >       ?                    @      �?              @        ������������������������       �                     @        @       A                   �Z@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        C       R       	          ����?\-��p�?"             M@       D       E                    @E@�<ݚ�?             B@        ������������������������       �                      @        F       Q       	          `ff�?@�0�!��?             A@       G       N                     Q@      �?             @@       H       M                    �? 	��p�?             =@        I       J                    a@r�q��?             (@       ������������������������       �                     @        K       L                   �l@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             1@        O       P                   pm@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        T       �       	          033�?�h��%�?�            `t@       U       r                    �?�
�@c�?�            �r@        V       g                   �c@v���EO�?0            �Q@       W       ^                   @E@     ��?              H@        X       ]                   �_@��
ц��?             *@       Y       \                   `[@�<ݚ�?             "@        Z       [                   �X@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        _       f                    �? >�֕�?            �A@       `       e       	          833�?$�q-�?             :@       a       b       	          ����?`2U0*��?             9@       ������������������������       �                     6@        c       d                   �j@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        h       k                    @I@�LQ�1	�?             7@        i       j                   �b@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        l       m                    m@�q�q�?             "@        ������������������������       �                     @        n       o                   �d@���Q��?             @        ������������������������       �                      @        p       q                   �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       �                   �g@@�沦~�?�            `l@       t       �                   �t@�/�z{�?�            @l@       u       �                    �? qP��B�?�            �j@        v       y                    �?��S�ۿ?             >@        w       x                   �`@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        z                          e@���7�?             6@       {       |                   �b@�����H�?             "@       ������������������������       �                     @        }       ~                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �       �                   `R@�x�V�?{             g@        �       �                    �?�����H�?             "@        �       �                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�|���?t             f@        ������������������������       �        '             Q@        �       �                   c@@3����?M             [@        �       �                   @[@`2U0*��?$             I@        ������������������������       �                     �?        �       �                   Hp@@�E�x�?#            �H@       ������������������������       �                     C@        �       �                   �p@�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        )             M@        �       �                    �?���!pc�?             &@        ������������������������       �                     @        �       �                   u@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �M@���>4��?             <@       �       �                   `U@ҳ�wY;�?             1@        ������������������������       �                     @        �       �                    �?�8��8��?             (@       �       �       	          ���@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@        �       �                   @o@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?F��_�?�             y@       �       �                    �?�I��Ǎ�?�             u@       �       �                   �V@�YnPB��?�            �p@        ������������������������       �                     �?        �       �                    Z@�!T���?�            �p@        ������������������������       �                    �F@        �       �                    \@��X��?�             l@        �       �                    `@���y4F�?             C@        �       �       
             �?���Q��?             $@        ������������������������       �                     @        �       �                   �Z@؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             �?@4և���?             <@        �       �                    @L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    `R@�nkK�?             7@       ������������������������       �                     4@        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   i@ rpa�?s            @g@        ������������������������       �        $             N@        �       �                   �\@�[|x��?O            �_@        �       �                   `_@�	j*D�?	             *@        ������������������������       �                     @        �       �                   �a@X�<ݚ�?             "@        �       �                   �`@      �?             @       �       �                   �k@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �Z@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ЮN
��?F            @\@        �       �                   �u@������?             .@       �       �                     H@8�Z$���?             *@        �       �                     F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     N@ףp=
�?
             $@       ������������������������       �                     @        �       �                    a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	          `ff�?@�E�x�?9            �X@       ������������������������       �                     K@        �       �       
             �?���7�?             F@        ������������������������       �                     "@        �       �                    c@ >�֕�?            �A@       ������������������������       �                     ?@        �       �                    q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?H�V�e��?+             Q@        �       �       	          033�?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �[@d�;lr�?'            �O@        �       �                   �Z@      �?              @        ������������������������       �                     @        �       �                   `Z@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?�C��2(�?"            �K@       �       �                   @e@�ݜ�?            �C@       �       �                   �b@�KM�]�?             C@       �       �                    n@�X�<ݺ?             B@       ������������������������       �                     4@        �       �                   �n@      �?	             0@        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        �             	             �?�P�*�?%             O@       �             	          ����?�q�q�?             B@       �                          0a@¦	^_�?             ?@       �       �                    �?      �?
             2@       �       �                   `]@�	j*D�?             *@        ������������������������       �                      @        �       �                    @K@"pc�
�?             &@       ������������������������       �                     @        �       �                    b@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     *@                                 �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                �^@$�q-�?             :@        ������������������������       �                     *@              
                   �?8�Z$���?	             *@              	                  p`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                 a@ףp=
�?             $@                                 @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  Ҙ
'�_�?��z���?�W�{��?P�� �?      �?     ��?z��y���?�0�0�?ާ�d��?C��6�S�?�Q����?
ףp=
�?              �?ffffff�?333333�?      �?              �?      �?      �?                      �?      �?      �?�؉�؉�?�;�;�?      �?                      �?ӛ���7�?d!Y�B�?      �?      �?      �?                      �?��y��y�?�a�a�?      �?                      �?�����?z�z��?��y��y�?�0�0�?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?        |���?|���?h/�����?&���^B�?      �?      �?      �?                      �?���Q��?)\���(�?UUUUUU�?UUUUUU�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?                      �?Y�B��?�Mozӛ�?�������?�������?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?              �?      �?              �?      �?              �?        F]t�E�?/�袋.�?      �?      �?              �?�������?�������?              �?      �?        �{a���?a����?�q�q�?9��8���?      �?        �������?ZZZZZZ�?      �?      �?�{a���?������?UUUUUU�?�������?              �?�������?333333�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?ǋ-����?��I� �?�ַC5�?�IA��U�?�
��V�?�ԓ�ۥ�?      �?      �?�؉�؉�?�;�;�?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ��+��+�?�A�A�?�؉�؉�?;�;��?���Q��?{�G�z�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        Nozӛ��?d!Y�B�?۶m۶m�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?q� 5��?����L�?H����?x�!���?��}A�?�}A_З?�������?�?      �?      �?      �?                      �?�.�袋�?F]t�E�?�q�q�?�q�q�?      �?              �?      �?              �?      �?              �?        ��5!({�?�	A����?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        ��.���?F]t�E�?      �?        ���Kh�?h/�����?���Q��?{�G�z�?              �?և���X�?9/���?      �?        ]t�E�?F]t�E�?              �?      �?              �?        F]t�E�?t�E]t�?      �?              �?      �?              �?      �?                      �?n۶m۶�?I�$I�$�?�������?�������?              �?UUUUUU�?UUUUUU�?]t�E�?F]t�E�?      �?                      �?      �?        F]t�E�?/�袋.�?�������?333333�?      �?                      �?              �?�z�G��?H�z�G�?�T�6|��?e�.y0��?= Y���?������?      �?        �%�N!�?P\[ ���?              �?%I�$I��?۶m۶m�?(������?6��P^C�?333333�?�������?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?        �$I�$I�?n۶m۶�?�������?�������?      �?                      �?d!Y�B�?�Mozӛ�?              �?UUUUUU�?UUUUUU�?              �?      �?        �n�ᆫ?Hy�G�?              �?EQEQ�?]�u]�u�?;�;��?vb'vb'�?              �?�q�q�?r�q��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?                      �?4��A�/�?m���M�?�?wwwwww�?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?      �?        9/���?և���X�?              �?F]t�E�?�.�袋�?              �?�A�A�?��+��+�?              �?      �?      �?              �?      �?        ZZZZZZ�?iiiiii�?333333�?�������?              �?      �?        �eY�eY�?��i��i�?      �?      �?      �?        333333�?�������?              �?      �?        F]t�E�?]t�E�?�i�i�?\��[���?(�����?�k(���?�q�q�?��8��8�?              �?      �?      �?      �?                      �?      �?              �?                      �?�Zk����?�RJ)���?UUUUUU�?UUUUUU�?��Zk���?�RJ)���?      �?      �?;�;��?vb'vb'�?      �?        F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?333333�?      �?                      �?;�;��?�؉�؉�?              �?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ܚihG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@@         ,                    �F@~jÚʞ�?<           ��@                                   �?�&KW���?}            �j@                                   �?����X�?-            �Q@                                  �E@䯦s#�?"            �J@                     
             �?��Q���?             D@                                  �D@ �Cc}�?             <@       ������������������������       �        	             0@                                   �?      �?             (@        	       
                   �[@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                  `m@�q�q�?	             (@                                 @^@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                      	             �?�	j*D�?	             *@                                  �?�����H�?             "@        ������������������������       �                     @                                  `i@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                  @]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@               #                    @�5?,R�?P             b@                                  �?PF��t<�?G            �_@        ������������������������       �                    �D@               "       
             �? �#�Ѵ�?/            �U@                !                   �b@����X�?             ,@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        '             R@        $       +                   �o@��.k���?	             1@       %       *                    �C@���!pc�?             &@       &       '                    e@���Q��?             @        ������������������������       �                      @        (       )       	          `ff�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        -       �       	          033�?L�9ͷ�?�            �@        .       c       
             �?r����w�?�            �u@        /       F                   `_@z[���?Z            `b@       0       C                   �o@�ɮ����?5            �V@       1       4       
             �?xdQ�m��?/            @T@        2       3                    @K@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        5       B                    @L@xL��N�?,            �R@        6       A                    �?�L���?            �B@       7       :                   `X@�C��2(�?            �@@        8       9                   �V@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ;       <                   �`@ 7���B�?             ;@       ������������������������       �                     3@        =       @                    �?      �?              @       >       ?                    @K@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �B@        D       E                    @O@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        G       R                    �?Dc}h��?%             L@        H       Q                    �?և���X�?
             ,@       I       P                    @O@���!pc�?             &@       J       O       	          ����?      �?              @       K       N                   `a@      �?             @        L       M                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        S       Z                    �?d}h���?             E@       T       U                    @L@���N8�?             5@       ������������������������       �        
             1@        V       Y       	          ����?      �?             @        W       X                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        [       ^                   �_@�ՙ/�?             5@        \       ]                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        _       `                   �c@؇���X�?             ,@       ������������������������       �                     $@        a       b                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        d       e       	          033��Mc��?}            @i@        ������������������������       �                     @        f       o                   @E@��2(&�?|            �h@        g       n                    �?      �?	             0@       h       k                    �?�eP*L��?             &@        i       j       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        l       m                   �b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        p       �                    �?�h�ഭ�?s            �f@        q       z                    �?������?            �F@        r       y                   �e@     ��?             0@       s       x                   Xv@      �?             (@       t       w                    �?ףp=
�?             $@       u       v                     K@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        {       |                    �?ܷ��?��?             =@        ������������������������       �                     @        }       ~                    �I@      �?             8@        ������������������������       �                     (@               �                    @J@      �?	             (@        �       �                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �c@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �g@���Z�?W             a@       �       �                    @L@г�wY;�?V             a@       ������������������������       �        8            @V@        �       �                   �^@dP-���?            �G@        ������������������������       �                     *@        �       �                   �_@�t����?             A@        ������������������������       �                     �?        �       �                     N@�C��2(�?            �@@        �       �                    �?�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                   pa@ �q�q�?             8@        ������������������������       �                     *@        �       �                   �s@�C��2(�?	             &@       ������������������������       �                     @        �       �                   �u@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�~f�7�?�            0v@       �       �                   �v@0G���ջ?�            @p@       �       �                    �H@0�`��!�?�            �o@        �       �                   @[@���B���?             :@        ������������������������       �                      @        �       �       	             �?      �?             8@        �       �                   @`@և���X�?             @        ������������������������       �                      @        �       �                    @H@z�G�z�?             @       �       �                    ]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        �       �       
             �?�u��?�            `l@        �       �       	             @��-�=��?            �C@        �       �                    �?���y4F�?             3@        �       �                    �?���!pc�?             &@        �       �       	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �N@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �Q@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    t@���e�?v            �g@       �       �                   �c@�E�����?q            �f@       �       �                    X@����?k            �e@        �       �                    �? ��WV�?             :@        ������������������������       �                     $@        �       �                    �?      �?             0@       ������������������������       �                     *@        �       �                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        _            @b@        �       �                   �d@      �?              @        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��C����?D            �W@        �       �                    �?�+e�X�?             9@        ������������������������       �                     @        �       �                   `c@�q�q�?             2@       �       �                   @q@$�q-�?             *@       ������������������������       �                     "@        �       �                   Xr@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?=��T�?2            �Q@       �       �       	           33@ҐϿ<��?*            �N@       �       �                    @N@�e�,��?)            �M@       �       �                   �q@���y4F�?             C@       �       �                   �e@6YE�t�?            �@@       �       �                   �`@      �?             @@        �       �                    �?������?
             1@        �       �       	          ���@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�8��8��?             (@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     .@        ������������������������       �                     �?        �       �       	          @33�?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    p@�G��l��?             5@       �       �                    @ҳ�wY;�?             1@       �       �                   �_@�q�q�?             (@       �       �                   �j@����X�?             @       �       �                    ]@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?z�G�z�?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �                           �?�q�q�?             "@       �       �       	          833@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B  g�����?L��/��?��~!V��?|d�S��?�$I�$I�?�m۶m��?�V�9�&�?�����?�������?333333�?۶m۶m�?%I�$I��?              �?      �?      �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?      �?        vb'vb'�?;�;��?�q�q�?�q�q�?      �?        �������?UUUUUU�?              �?      �?              �?      �?      �?                      �?              �?�q�q�?�q�q�?�������?�@ �?      �?        �/����?�}A_Ч?�m۶m��?�$I�$I�?              �?      �?              �?        �?�������?F]t�E�?t�E]t�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?t�E]t�?F]t�E�?h�5#�?0�甹��?�E�_���?��(W�?�Q�Q�?]��\���?X�<ݚ�?�5?,R�?�$I�$I�?�m۶m��?      �?                      �?L�Ϻ��?>�S��?L�Ϻ��?}���g�?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?        h/�����?	�%����?              �?      �?      �?�$I�$I�?۶m۶m�?              �?      �?                      �?              �?              �?�������?333333�?              �?      �?        ۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?              �?                      �?۶m۶m�?I�$I�$�?�a�a�?��y��y�?              �?      �?      �?      �?      �?      �?                      �?              �?�a�a�?�<��<��?۶m۶m�?�$I�$I�?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?5r���?+�7����?              �?��.���?t�E]t�?      �?      �?t�E]t�?]t�E�?�������?�������?      �?                      �?�������?UUUUUU�?      �?                      �?              �?-�-��?�~�~�?wwwwww�?�?      �?      �?      �?      �?�������?�������?UUUUUU�?�������?      �?                      �?              �?      �?              �?        ��=���?a���{�?      �?              �?      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?      �?                      �?�J���?T{N���?�?�?      �?        �����F�?W�+�ɵ?      �?        <<<<<<�?�?              �?]t�E�?F]t�E�?9��8���?�q�q�?              �?      �?        �������?UUUUUU�?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?                      �?8&yȎ��?r��M\��?�؉�؉�?vb'vb'�?'���H�?.Wr{�?ى�؉��?��؉���?      �?              �?      �?۶m۶m�?�$I�$I�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?{��U���?tSRb�?�A�A�?}˷|˷�?(������?6��P^C�?t�E]t�?F]t�E�?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?                      �?AL� &W�?����F}�?l�l��?P��O���?�}A_�w?�}A_��?;�;��?O��N���?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?        ��%N��?#�X��?R���Q�?���Q��?      �?        UUUUUU�?UUUUUU�?�؉�؉�?;�;��?      �?              �?      �?              �?      �?                      �?�������?�:��:��?mާ�d�?������?_[4��?�pR���?(������?6��P^C�?e�M6�d�?'�l��&�?      �?      �?�?xxxxxx�?333333�?�������?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        333333�?�������?      �?                      �?1�0��?��y��y�?�������?�������?�������?�������?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���+hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�D         �       
             �?T �����?N           ��@              -                    �?��U�E�?H           �@               &                    �?      �?1            �S@              %       	          033@�U���?%             O@                                 @]@~|z����?             �J@                                   �?�8��8��?             (@                                  �?z�G�z�?             @        ������������������������       �                      @        	       
                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                  @b@v�2t5�?            �D@                     
             �?������?             ;@        ������������������������       �                      @                                   �?z�G�z�?             9@                                 �V@      �?
             4@        ������������������������       �                      @                                   �?r�q��?	             2@                     	          ����?��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@                                  @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               $                    �?����X�?             ,@              #       	          ����?�q�q�?
             (@              "                    �?���Q��?             $@              !       	          @33�?�q�q�?             @                                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        '       ,                   0e@      �?             0@       (       )                    �?��S�ۿ?             .@        ������������������������       �                     @        *       +                   �h@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        .       k                    �?������?           �z@       /       \                   �b@�v�\�?�             s@       0       Y                    �R@����,��?�            �q@       1       2       	            �?H��2�?�            pq@        ������������������������       �        )             M@        3       4                    �?0�%�J�?�            �k@        ������������������������       �                    �B@        5       R                    @M@���.�6�?t             g@       6       7                   �U@̹�"���?E            �[@        ������������������������       �                     �?        8       I                    @L@�C��2(�?D            �[@       9       B                    �?�X�<ݺ?6            �V@       :       =                     E@�i�y�?)            �O@        ;       <                     D@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        >       A                    �?0�)AU��?%            �L@        ?       @                   hq@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                    �G@        C       H                   �_@�����H�?             ;@        D       G       	             @���Q��?             @       E       F                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             6@        J       M       	          ����?      �?             4@        K       L                    X@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        N       Q                   �i@$�q-�?	             *@        O       P                    ^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        S       X                   �`@ �й���?/            @R@        T       W       	             �? ��WV�?             :@        U       V                    �O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     �G@        Z       [                   �b@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ]       ^       	          833�?���!pc�?             6@        ������������������������       �                     @        _       f                    �?�q�q�?             2@        `       a                   pd@�eP*L��?             &@        ������������������������       �                     @        b       c                   �e@؇���X�?             @        ������������������������       �                     @        d       e                   @Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        g       h                   �`@؇���X�?             @        ������������������������       �                     @        i       j                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       }                   a@��
��X�?O            @_@        m       |                    �?     p�?$             P@       n       q                    �E@�Ra����?             F@        o       p                    �C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        r       y                   �s@��p\�?            �D@       s       x                   �\@�7��?            �C@        t       w                    �?"pc�
�?             &@        u       v       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     <@        z       {                    �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        ~       �                    �?x>ԛ/��?+            �N@               �                   q@�q�q�?             8@       �       �                    @L@R���Q�?             4@        ������������������������       �                     &@        �       �                    �N@�q�q�?             "@       �       �       	          ���@���Q��?             @       �       �                   Pc@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @E@4�B��?            �B@        �       �                    ]@����X�?             @        ������������������������       �                     @        �       �                   �l@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�������?             >@       �       �                    �?��s����?             5@       �       �                    �?      �?             0@       �       �                    �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �       	            �?      �?             @        ������������������������       �                     �?        �       �                   f@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @M@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�|�LH��?           �y@       �       �                    �?>��i3�?�            0u@        �       �                   �u@���g�?D            �Y@       �       �                    �?�q�q�?@             X@        �       �                    k@���@M^�?             ?@        ������������������������       �                     @        �       �                    �L@�q�����?             9@       �       �                     D@     ��?	             0@        ������������������������       �                     @        �       �                   `t@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �c@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   @^@@i��M��?.            @P@        �       �                   `T@@4և���?             ,@        �       �                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �X@x�K��?!            �I@        ������������������������       �                     @        �       �                    `@"Ae���?            �G@        �       �       	             �?���!pc�?             &@        �       �                    m@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �P@�<ݚ�?             B@       �       �                   `a@6YE�t�?            �@@        ������������������������       �        	             (@        �       �                   pf@���N8�?             5@       �       �       	             �?�S����?             3@       �       �       	             �?�θ�?	             *@       �       �                    @K@r�q��?             (@        ������������������������       �                     @        �       �                   �c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?Xc!J�ƴ?�            �m@        �       �                    �?4?,R��?             B@       �       �                    @     ��?             @@       �       �                     H@�>����?             ;@        ������������������������       �                     @        �       �                    �?ףp=
�?             4@        ������������������������       �                     @        �       �                   �]@�t����?             1@        �       �                    j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �d@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        �       �       	          ����?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    I@�(\����?�             i@        �       �                   pf@�q�q�?             "@       �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    @ bj�p8�?z            �g@       ������������������������       �        p            �e@        �       �                   �c@      �?
             0@        ������������������������       �                      @        �       �                   0i@      �?              @        ������������������������       �                     @        �       �                   �a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �]@��(@��?*            �Q@        �       �                    `P@�<ݚ�?	             2@       �       �                   �l@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     @        �                          �M@����3��?!             J@       �       �                   `R@      �?             B@        ������������������������       �                     @        �       �                   `]@ףp=
�?             >@        ������������������������       �                     �?        �                          �? 	��p�?             =@       �                          �? 7���B�?             ;@                                  �?ףp=
�?             $@                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@                                 �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	      
                   �?      �?             0@        ������������������������       �                     @                                 �?�θ�?	             *@                               �b@�z�G��?             $@                                �?      �?              @        ������������������������       �                     @                    	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KMKK��hb�B0  ��G��G�?�\�\�?���/u��? �"�?      �?      �?�9�s��?c�1��?��sHM0�?�	�[���?UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?��+Q��?�ڕ�]��?B{	�%��?{	�%���?              �?�������?�������?      �?      �?              �?�������?UUUUUU�?�������?�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?�������?333333�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?              �?              �?      �?      �?�������?�?      �?        �q�q�?�q�q�?              �?      �?                      �?r��U�?}������?�������?�������?Zas �
�?����RO�?X`��?�~�駟�?              �?�ͫ?~/C~/C�?              �?Y�B��?���7���?镱��^�?C�I .��?      �?        F]t�E�?]t�E�?�q�q�?��8��8�?AA�?�������?UUUUUU�?�������?              �?      �?        p�}��?��Gp�?�������?�������?              �?      �?                      �?�q�q�?�q�q�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?�$I�$I�?۶m۶m�?              �?      �?        ;�;��?�؉�؉�?      �?      �?      �?                      �?              �?����?����Ǐ�?;�;��?O��N���?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?333333�?�������?              �?      �?        t�E]t�?F]t�E�?              �?UUUUUU�?UUUUUU�?]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?�� �rh�?����K�?      �?     ��?]t�E�?]t�E]�?UUUUUU�?UUUUUU�?              �?      �?        ��+Q��?�]�ڕ��?�A�A�?��[��[�?F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?              �?      �?      �?              �?      �?                      �?�K�`m�?;ڼOq��?�������?�������?333333�?333333�?      �?        UUUUUU�?UUUUUU�?�������?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?              �?                      �?L�Ϻ��?�Y7�"��?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?�������?�������?�a�a�?z��y���?      �?      �?F]t�E�?]t�E�?      �?                      �?333333�?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?         U8����?������?�{���G�?�.�	��?^�	���?C����?�������?�������?�c�1��?�s�9��?              �?���Q��?�p=
ף�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?      �?        �Z��Z��?�J��J��?n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?        ssssss�?�?              �?�w6�;�?W�+���?t�E]t�?F]t�E�?      �?      �?      �?                      �?              �?9��8���?�q�q�?'�l��&�?e�M6�d�?      �?        �a�a�?��y��y�?(������?^Cy�5�?ى�؉��?�؉�؉�?�������?UUUUUU�?      �?        333333�?�������?      �?                      �?              �?      �?                      �?              �?      �?        �؊���?�pR�履?�8��8��?r�q��?      �?      �?�Kh/��?h/�����?      �?        �������?�������?      �?        <<<<<<�?�?      �?      �?              �?      �?        �������?�?      �?                      �?�������?333333�?              �?      �?              �?        333333�?�������?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?S�K8��?:kP<�q�?      �?              �?      �?      �?              �?      �?      �?        333333�?�������?              �?      �?        ����?��+��+�?�q�q�?9��8���?�?�������?              �?      �?              �?        ��N��N�?'vb'vb�?      �?      �?              �?�������?�������?              �?������?�{a���?	�%����?h/�����?�������?�������?      �?      �?              �?      �?              �?              �?              �?      �?      �?                      �?      �?      �?      �?        �؉�؉�?ى�؉��?333333�?ffffff�?      �?      �?              �?      �?      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ4��chG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�C         �       
             �?�>�Ļ`�?N           ��@                                  �F@>�H�{�?T           ��@                                  �c@@i��M��?+            @P@                                  �?�T|n�q�?            �E@              
                   �j@      �?             @@                                  Pb@      �?             0@       ������������������������       �        	             ,@               	                    Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@                                   @�eP*L��?             &@                                 �p@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                   @C@���|���?             6@                     
             �?�q�q�?             (@        ������������������������       �                     @                                  �f@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@               )                   f@��|��?)           @}@               &                   �c@@A��q�?P            �`@                                 `\@ qP��B�?M             `@                                  ``@�KM�]�?             3@       ������������������������       �                     1@        ������������������������       �                      @               %                    �?����r�?A            �[@              $       
             �?����e��?'            �P@                #                    �?ףp=
�?             $@        !       "                   �T@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        "             L@        ������������������������       �                     F@        '       (                   0d@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        *       S                    �?x�)Z	e�?�            �t@        +       H                    �?T�7�s��?(            �L@       ,       =                   �a@������?            �D@       -       0                    �?      �?             4@        .       /       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        1       <                   �`@���Q��?
             .@       2       9                    s@      �?             (@       3       4                   @[@����X�?             @        ������������������������       �                     �?        5       8                   �q@r�q��?             @        6       7                   l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        :       ;       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        >       E                   u@�����?             5@       ?       D       	          ����?�}�+r��?             3@       @       C                   pl@@4և���?             ,@        A       B                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     @        F       G                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       J                   `X@     ��?             0@        ������������������������       �                     �?        K       R                   �`@�r����?             .@       L       Q                    �?����X�?             @        M       N       	             �?�q�q�?             @        ������������������������       �                     �?        O       P                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        T       �                   �a@8zw"׷�?�            @q@       U       ~                   Pz@�X�<ݺ?�             k@       V       o                   ``@� Λ��?�            �j@        W       n       	          ����?��O���?9            @U@       X       Y       	          ����?:	��ʵ�?             �F@        ������������������������       �                     1@        Z       m                    �P@����X�?             <@       [       h                    �O@�q�q�?             8@       \       g                    �?���y4F�?             3@       ]       f                     M@r�q��?             2@        ^       _                   @i@      �?             @        ������������������������       �                     �?        `       e                    @L@���Q��?             @       a       d                    �?      �?             @        b       c                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        i       j       	             �?z�G�z�?             @        ������������������������       �                     @        k       l                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     D@        p       w       	          ����? qP��B�?P             `@        q       r                    �?ףp=
�?             4@        ������������������������       �                     (@        s       v                   �\@      �?              @        t       u                     N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        x       y                    �?��wڝ�?D            @[@       ������������������������       �        -            �S@        z       }                   `\@�g�y��?             ?@        {       |                     R@ףp=
�?	             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     5@               �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?&             N@        �       �                    �?��2(&�?             6@       �       �                   �a@      �?             (@       �       �                    �?      �?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                     I@D�n�3�?             C@        ������������������������       �                     @        �       �                   �b@�q�q�?            �@@        �       �                   b@��.k���?
             1@        �       �                   �a@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �a@�<ݚ�?             "@       �       �                    �K@      �?              @        �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �L@     ��?
             0@       ������������������������       �                     $@        �       �       	          ����?      �?             @       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �O@z�G�z�?�            x@        �       �                    @M@��>4և�?!             L@       �       �                   �`@H�V�e��?             A@       �       �       	          ����?��� ��?             ?@        �       �                   �W@�q�q�?             (@        ������������������������       �                     @        �       �                    �?      �?              @        �       �       	          �����q�q�?             @        ������������������������       �                     �?        �       �                   Pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �F@���Q��?             @       �       �                    @D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             3@        ������������������������       �                     @        �       �       	          `ff�?�X����?             6@       �       �                    �?     ��?	             0@       �       �                   �c@�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                    a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @L@0�5��?�            �t@       �       �       	             �?j��pX�?�             o@       �       �                    �?�G���?�            �k@        �       �                    �?>a�����?!            �I@       �       �                    �? �#�Ѵ�?            �E@        ������������������������       �                     (@        �       �                   �l@`Jj��?             ?@        ������������������������       �        	             0@        �       �       	          ����?�r����?             .@       �       �                   `\@8�Z$���?
             *@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    @G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @n@��$����?v            �e@       ������������������������       �        I            @Z@        �       �                    �?�����?-            �P@        ������������������������       �                     $@        �       �                   0c@�}�+r��?&            �L@        �       �                   �\@��2(&�?             6@        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                    �A@        �       �                   �u@�+e�X�?             9@       �       �       	          ����?�㙢�c�?             7@        �       �                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   hq@�KM�]�?             3@       �       �                   �c@��S�ۿ?             .@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�w���?2            @T@        �       �                    �N@��2(&�?             6@        �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     .@        �                          �?Ɣ��Hr�?%            �M@       �       �                   �h@�5��
J�?             G@        ������������������������       �                     *@        �                          @�q�q�?            �@@       �       �                   �i@      �?             <@        ������������������������       �                      @        �       �                   0c@���B���?             :@       ������������������������       �                     2@        �       �                   �k@      �?              @        ������������������������       �                     �?        �                          �?����X�?             @                                 �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                    	          @33�?z�G�z�?             @        ������������������������       �                      @                                �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        	                        �_@$�q-�?
             *@        
                         @N@z�G�z�?             @        ������������������������       �                     @                                 \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  Qm4��?X��;�?�m�u���?��"���?�J��J��?�Z��Z��?6eMYS��?���)k��?      �?      �?      �?      �?              �?      �?      �?              �?      �?                      �?t�E]t�?]t�E�?      �?      �?      �?                      �?              �?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?      �?              �?        � � �?˷|˷|�?t��:W�?��)F�?�}A_З?��}A�?(�����?�k(���?              �?      �?        ��)A��?�oX����?|���?�>����?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?UUUUUU�?�������?      �?                      �?O}Q����?��kD�
�?�}��?p�}��?��+Q��?�v%jW��?      �?      �?�������?�������?      �?                      �?�������?333333�?      �?      �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?                      �?              �?�a�a�?=��<���?(�����?�5��P�?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?              �?      �?              �?      �?              �?�������?�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?        ?���(�?;0�̵�?�q�q�?��8��8�?7��XQ�?�L�w�Z�?�?�������?l�l��?��O��O�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?(������?6��P^C�?UUUUUU�?�������?      �?      �?      �?        �������?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?      �?        �������?�������?      �?              �?      �?              �?      �?                      �?              �?�}A_З?��}A�?�������?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�,�M�ɂ?N��ش�?              �?�B!��?��{���?�������?�������?              �?      �?                      �?      �?      �?      �?                      �?�������?�������?t�E]t�?��.���?      �?      �?      �?      �?              �?      �?      �?      �?              �?      �?              �?      �?                      �?              �?l(�����?(������?              �?UUUUUU�?UUUUUU�?�������?�?      �?      �?      �?                      �?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?              �?      �?      �?              �?      �?      �?      �?      �?                      �?              �?�������?�������?I�$I�$�?۶m۶m�?ZZZZZZ�?iiiiii�?�B!��?�{����?UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �E]t��?]t�E]�?      �?      �?�������?�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�{Y%P��?�j���?�9�s��?�1�c��?_�T
�k�?ʰZoA�?�������?�?�/����?�}A_Ч?      �?        ���{��?�B!��?      �?        �������?�?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?      �?              �?      �?        �w�q�?w�qGܑ?      �?        g��1��?���@��?      �?        �5��P�?(�����?��.���?t�E]t�?              �?      �?              �?        R���Q�?���Q��?�7��Mo�?d!Y�B�?      �?      �?              �?      �?        �k(���?(�����?�������?�?�������?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?              �?��Hx��?�n���?��.���?t�E]t�?�$I�$I�?۶m۶m�?              �?      �?              �?        ��c+���?#h8����?�,d!Y�?�Mozӛ�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?��؉���?ى�؉��?      �?              �?      �?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?�؉�؉�?�������?�������?              �?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���=hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK�h��B�<         �                    �?z�ГPo�?D           ��@              c       
             �?�8<L��?C           �@              `                    �R@�^'�ë�?�            @x@                     	          833�?`�,"��?�            �w@        ������������������������       �        .             T@                                   �?�/oD�?�            �r@                                   �?v�X��?              F@               	                    @K@�G�z��?             4@        ������������������������       �                     @        
              	          ����?8�Z$���?	             *@                                   �O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@                      	          ����?r�q��?             8@                                   �?      �?             @                     	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                    Q@ףp=
�?             4@                     	          033�?�}�+r��?             3@       ������������������������       �                     1@                      	          ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               !       	          ����?�}�}CS�?�            0p@                                    �?����X�?             @                                 �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        "       ]                   �z@�[|x��?�            �o@       #       \                   �c@j��pX�?�             o@       $       [                   �r@��q���?�            �n@       %       X                   `r@$�q-�?�             j@       &       Q                   Pb@�/a��I�?�            �i@       '       P                    �?�IєX�?}            `g@       (       C       	          ����?pOW�1J�?Y            �`@        )       8       	          033�?PN��T'�?!             K@       *       /       	          ����?�}�+r��?             C@        +       .                    �?z�G�z�?             @       ,       -                   �_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        0       1                    �?Pa�	�?            �@@       ������������������������       �                     <@        2       7       	          033�?z�G�z�?             @       3       6                   �j@      �?             @       4       5                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        9       :                   �]@      �?
             0@        ������������������������       �                     @        ;       <                    �?�eP*L��?             &@        ������������������������       �                      @        =       @                    �K@X�<ݚ�?             "@       >       ?                    @G@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        A       B                   @`@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        D       I       
             �?x�G�z�?8             T@        E       H       	          ��� @��S�ۿ?             .@        F       G                    Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             (@        J       K       	          033@��ɉ�?-            @P@       ������������������������       �                     �F@        L       O                   �_@ףp=
�?             4@        M       N       	          ���@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             .@        ������������������������       �        $            �J@        R       U                    @L@r�q��?	             2@       S       T                   �Z@@4և���?             ,@        ������������������������       �                     �?        ������������������������       �                     *@        V       W                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        Y       Z                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �C@        ������������������������       �                     �?        ^       _                   @X@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        a       b       
             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        d       �       	          ����?�lhM��?O            �_@       e       l                    �?����X�?/            @S@        f       k                   xt@�����H�?
             2@       g       h                    s@�IєX�?	             1@       ������������������������       �                     ,@        i       j                    e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        m       �                    �?L
�q��?%            �M@       n       y                    �?R�}e�.�?!             J@       o       p                   �b@�����H�?             B@       ������������������������       �                     5@        q       x                    �K@������?	             .@       r       u                    �?���|���?             &@        s       t                   �f@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        v       w                   q@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        z                          �b@      �?
             0@        {       ~                    �?z�G�z�?             @        |       }                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?"pc�
�?             &@        �       �                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @`@�����H�?             "@        ������������������������       �                     @        �       �                    a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �p@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   ``@H.�!���?              I@        �       �                    @M@�nkK�?             7@       �       �                     L@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?��}*_��?             ;@        �       �                   �V@�θ�?	             *@        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �        	             ,@        �       �       	          ����?F��Y���?           0y@       �       �                   �X@��3E��?�            pq@        �       �       
             �?�q�q�?
             2@       ������������������������       �                     (@        ������������������������       �                     @        �       �                    @L@�N��D�?�            Pp@       �       �                    I@�7A��?�             i@        �       �                   @^@z�G�z�?             @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?�Q �?�            �h@        �       �                    �?*;L]n�?             >@       �       �                   `a@$��m��?             :@       �       �                   �n@��s����?             5@       ������������������������       �                     (@        �       �                    �?X�<ݚ�?             "@       �       �                   �a@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        p            �d@        �       �                   pk@d��0u��?"             N@        �       �       	          ����?���Q��?             9@        �       �                    @M@8�Z$���?             *@        ������������������������       �                     @        �       �                    X@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       	            �?�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        �       �                   �c@z�G�z�?            �A@       �       �                   �m@ �Cc}�?             <@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     6@        �       �       
             �?և���X�?             @       �       �                   8p@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �_@�g�y��?L             _@        �       �                    �?      �?             B@        �       �                   �n@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   `_@\-��p�?             =@        �       �                   �Z@���!pc�?             &@        ������������������������       �                     @        �       �                   �j@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�X�<ݺ?             2@        �       �                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             .@        �       �                   �d@      �?5             V@        ������������������������       �                     $@        �       �                   �o@^Gث3��?/            �S@       �       �       	          ���@      �?              L@       �       �                    �?��<D�m�?            �H@        ������������������������       �                     ,@        �       �       	          ��� @�#-���?            �A@       �       �                   @h@�IєX�?             A@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �^@ 7���B�?             ;@        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                    @J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             1@        ������������������������       �                     �?        �       �                   @n@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                   0r@���!pc�?             6@       �       �                   0q@�S����?             3@        ������������������������       �                     "@        �       �                    �?�z�G��?             $@        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  1�i�M��?��<Y �?�_G{X�?�:.�i�?���Id�?=�L�v��?l�s-Df�?��Qz7��?              �?�옥��?�ę֞��?颋.���?�.�袋�?�������?�������?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?(�����?�5��P�?              �?      �?      �?      �?                      �?      �?        ^��d޵�?��e3D��?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?        EQEQ�?]�u]�u�?�1�c��?�9�s��?T	9?��?���X��?;�;��?�؉�؉�?|��{�?ѽ݋��?�?�?~5&��?=P9��_�?h/�����?&���^B�?(�����?�5��P�?�������?�������?      �?      �?              �?      �?                      �?|���?|���?              �?�������?�������?      �?      �?      �?      �?      �?                      �?              �?              �?      �?      �?              �?t�E]t�?]t�E�?      �?        �q�q�?r�q��?�������?�������?      �?                      �?      �?      �?      �?                      �?333333�?�������?�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �? �����??�?��?              �?�������?�������?�������?333333�?      �?                      �?              �?              �?UUUUUU�?�������?�$I�$I�?n۶m۶�?      �?                      �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?      �?                      �?�������?333333�?      �?                      �?(
�B��?����z��?�m۶m��?�$I�$I�?�q�q�?�q�q�?�?�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?��V'�?�pR���?'vb'vb�?�;�;�?�q�q�?�q�q�?      �?        wwwwww�?�?]t�E]�?F]t�E�?�������?333333�?              �?      �?        �������?UUUUUU�?              �?      �?              �?              �?      �?�������?�������?      �?      �?              �?      �?              �?        F]t�E�?/�袋.�?      �?      �?      �?                      �?�q�q�?�q�q�?              �?�������?�������?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?        )\���(�?�(\����?d!Y�B�?�Mozӛ�?F]t�E�?]t�E�?              �?      �?                      �?B{	�%��?_B{	�%�?ى�؉��?�؉�؉�?              �?      �?                      �?~����/�?����?'�h��&�?f�]v�e�?UUUUUU�?UUUUUU�?              �?      �?        �~�u�7�?�2)^ �?nZq�$K�?�,u�ئ�?�������?�������?      �?      �?      �?                      �?              �?x9/���??4և���?""""""�?�������?�N��N��?vb'vb'�?z��y���?�a�a�?      �?        r�q��?�q�q�?�m۶m��?�$I�$I�?              �?      �?                      �?              �?              �?      �?        DDDDDD�?wwwwww�?�������?333333�?;�;��?;�;��?              �?�$I�$I�?�m۶m��?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?%I�$I��?۶m۶m�?      �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?                      �?              �?�B!��?��{���?      �?      �?�m۶m��?�$I�$I�?      �?                      �?�{a���?a����?t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?                      �?�q�q�?��8��8�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?i�i��?�-��-��?      �?      �?��S�r
�?և���X�?      �?        �A�A�?_�_�?�?�?۶m۶m�?�$I�$I�?      �?                      �?	�%����?h/�����?�������?�������?      �?              �?      �?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?        t�E]t�?F]t�E�?^Cy�5�?(������?              �?333333�?ffffff�?              �?      �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ--7BhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@@         *                    _@>���i��?F           ��@                      
             �?B�xX�?m            `d@              
                    �J@��u}���?Q            �]@               	       
             �?�S����?             C@                                   �?�eP*L��?             &@        ������������������������       �                     @                                   @J@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ;@                                   �Q@ 7���B�?8            @T@                                  �? ���J��?5            �S@       ������������������������       �        $             K@                                   @O@�8��8��?             8@       ������������������������       �                     1@                      	          ����?����X�?             @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                      
             �?�q�q�?             @        ������������������������       �                     �?                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               )                   0f@�X���?             F@                                 `]@������?            �D@        ������������������������       �                     $@               "                   �_@���@M^�?             ?@                                   �?r�q��?             (@        ������������������������       �                      @                !                     P@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        #       (                    �?�\��N��?             3@       $       %                    �?r�q��?             (@       ������������������������       �                      @        &       '       	             �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        +       �       	             �?������?�           ��@       ,       g                    �L@��;q�?�            �x@       -       <                    �F@�;n��?�            @s@        .       3       
             �?,mG����?U             `@        /       0                    �?      �?             0@        ������������������������       �                     @        1       2                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        4       ;                   `\@ T���v�?I            @\@        5       6                   pb@�S����?             3@        ������������������������       �                     @        7       :                    �?�θ�?	             *@        8       9                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        <            �W@        =       ^                    �?�0ϔ'6�?m            `f@       >       K       
             �?z���=��?^            @c@        ?       D                    �?���@M^�?             ?@        @       A       	          ����?      �?	             0@       ������������������������       �                     *@        B       C                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        E       F                    �?�q�q�?	             .@        ������������������������       �                     @        G       J                    �?X�<ݚ�?             "@       H       I                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        L       M                   �l@��sK�z�?L            �^@       ������������������������       �        (             Q@        N       U                    ]@X�;�^o�?$            �K@        O       T                    �?�q�q�?             .@       P       Q                   �b@�eP*L��?             &@        ������������������������       �                     @        R       S                   o@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        V       ]                   @g@P���Q�?             D@       W       X                   pd@ ���J��?            �C@       ������������������������       �                     ?@        Y       \                    �?      �?              @        Z       [                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        _       f       
             �?� �	��?             9@       `       a                   �`@      �?
             0@        ������������������������       �                     @        b       c                     H@�<ݚ�?             "@        ������������������������       �                     �?        d       e                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        h       �                    �?և���X�?7             U@       i       v       
             �?��y�:�?+            �P@        j       u                    �Q@      �?             8@       k       p                    �?�\��N��?
             3@        l       o                   �l@�q�q�?             (@       m       n                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        q       r                    �?����X�?             @        ������������������������       �                     @        s       t                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        w       �                    �?�T|n�q�?            �E@        x       }                    �?��
ц��?
             *@        y       |                   �u@����X�?             @       z       {                   f@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ~                          �h@r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �s@(;L]n�?             >@       ������������������������       �                     <@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?@�0�!��?             1@       ������������������������       �                     (@        �       �                   0`@���Q��?             @       �       �                    �O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?@b�?�            �v@       �       �                    �?�����?�            �o@        �       �                    �?R�}e�.�?             J@       �       �                   0e@��k=.��?            �G@       �       �       
             �?��2(&�?             F@       �       �                    �Q@�KM�]�?             C@       �       �                    �?�L���?            �B@        �       �                    �M@P���Q�?
             4@        �       �                    �?z�G�z�?             @       �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        �       �                   �`@�t����?             1@        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        �       �       	          ����?z�G�z�?             @        �       �                   `Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �a@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   P`@P���Q�?y             i@        �       �                    �?�̨�`<�?4            @U@        �       �                   �\@��
ц��?             *@        ������������������������       �                     @        �       �                    @I@���Q��?             $@        ������������������������       �                      @        �       �                   �r@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �? �q�q�?-             R@       �       �                   Pi@P����?#            �M@        �       �                   �h@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                    �E@        �       �       
             �?8�Z$���?
             *@        ������������������������       �                     @        �       �                   �q@�<ݚ�?             "@       �       �       	             �?      �?             @        ������������������������       �                     �?        �       �       	             @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    q@@���a��?E            �\@       ������������������������       �        +            �P@        �       �                    �?@��8��?             H@        ������������������������       �                     0@        �       �                   0q@      �?             @@        �       �                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     >@        �       �                    �?�f��`��?I            �[@       �       �       	          ���@�Pf����??            �W@       �       �                   �`@=&C��?5            �T@        �       �                   @Y@�<ݚ�?             2@        ������������������������       �                      @        �       �                   `^@      �?             0@        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   r@�θ�?(            @P@       �       �                   0o@���3�E�?!             J@       �       �                    @P@�MI8d�?            �B@       �       �                   �g@�t����?             A@        �       �       
             �?և���X�?             @        ������������������������       �                     @        �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �m@ 7���B�?             ;@       ������������������������       �                     2@        �       �                    �?�����H�?             "@       ������������������������       �                     @        �       �                    n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          `ff�?���Q��?	             .@       �       �                   `q@�q�q�?             "@        ������������������������       �                     @        �       �       
             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        �       �                   �p@r�q��?
             (@       �       �       	          ���
@�C��2(�?	             &@       ������������������������       �                     @        �       �       	          `ff@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?
             0@        ������������������������       �                     �?        �                           �?��S�ۿ?	             .@        �       �                   �h@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �t�bh�h)h,K ��h.��R�(KMKK��hb�B  �Q��Q��?W�W��?��\w���?��(��I�?�\�\�?�o��o��?^Cy�5�?(������?t�E]t�?]t�E�?      �?              �?      �?              �?      �?                      �?h/�����?	�%����?�A�A�?��-��-�?              �?UUUUUU�?UUUUUU�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�E]t��?]t�E�?��+Q��?�v%jW��?              �?�c�1��?�s�9��?UUUUUU�?�������?              �?�������?�������?              �?      �?        y�5���?�5��P�?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �5[g�?-�I��1�?9/����?�Cc}h�?!��O���?{����1�?QW�uE�?uE]QWԵ?      �?      �?      �?        �q�q�?�q�q�?              �?      �?        6h�e�&�?4��A�/�?(������?^Cy�5�?      �?        ى�؉��?�؉�؉�?      �?      �?      �?                      �?      �?              �?        ��z�b��?�Fu��?�cj`��?
qV~B��?�c�1��?�s�9��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?        �q�q�?r�q��?      �?      �?      �?                      �?              �?.����-�?#6�a#�?      �?        �־a��?J��yJ�?UUUUUU�?UUUUUU�?t�E]t�?]t�E�?      �?        �$I�$I�?�m۶m��?              �?      �?              �?        ffffff�?�������?��-��-�?�A�A�?      �?              �?      �?      �?      �?              �?      �?              �?                      �?)\���(�?�Q����?      �?      �?              �?�q�q�?9��8���?      �?              �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?�@��~�?~5&��?      �?      �?�5��P�?y�5���?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?���)k��?6eMYS��?�;�;�?�؉�؉�?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?              �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�?      �?              �?      �?              �?      �?        �������?ZZZZZZ�?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        vK�B#��?#-@/w��?�a�a�?=��<���?�;�;�?'vb'vb�?br1���?g���Q��?t�E]t�?��.���?(�����?�k(���?L�Ϻ��?}���g�?�������?ffffff�?�������?�������?      �?      �?      �?                      �?              �?              �?�?<<<<<<�?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?              �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �������?ffffff�?�?�������?�؉�؉�?�;�;�?              �?333333�?�������?      �?              �?      �?      �?                      �?UUUUUU�?�������?'u_[�?�V'u�?      �?      �?              �?      �?                      �?;�;��?;�;��?              �?�q�q�?9��8���?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?���ρ?�uI�ø�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?      �?                      �?              �?�5'���?�蕱���?�-q����?a�+F�?�%���?�����\�?�q�q�?9��8���?      �?              �?      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?ى�؉��?�؉�؉�?O��N���?b'vb'v�?��L���?L�Ϻ��?<<<<<<�?�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?        	�%����?h/�����?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        UUUUUU�?�������?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?      �?              �?      �?      �?        �?�������?�������?�������?      �?                      �?              �?�t�bub�
+     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJCM�,hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK煔h��B�9         �                    �?�7i���?A           ��@              A                   �`@$aA3yl�?;           �~@                                  �?��� ��?�            �r@                                   �N@��
ц��?             :@                                 �`@D�n�3�?             3@                                 �X@"pc�
�?             &@        ������������������������       �                     �?               	                    �?ףp=
�?             $@       ������������������������       �                     @        
                          @_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                      	             �?      �?              @        ������������������������       �                      @        ������������������������       �                     @                                  �R@؇���X�?             @        ������������������������       �                     @                                  @_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               *       	            �?ДX��?�             q@               )                    �?������?*            �R@              $                   �a@ڡR����?            �H@              #       	          833�?p9W��S�?             C@                                  Z@      �?             B@                                   �?      �?             0@                                  U@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @               "                   �[@P���Q�?             4@                !                   0j@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                      @        %       &       
             �?"pc�
�?             &@        ������������������������       �                     �?        '       (                    Z@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     :@        +       6                    �?���ؑ�?}            �h@        ,       1       	          ����?      �?             @@        -       .                   �_@���!pc�?             &@        ������������������������       �                     @        /       0       
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        2       5       
             �?���N8�?             5@        3       4                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     3@        7       >                   @X@�'���8�?h            �d@        8       =                   �`@؇���X�?
             ,@        9       :                    �K@�q�q�?             @        ������������������������       �                     @        ;       <                   Pl@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ?       @                    �R@ 1�P<Ě?^            �b@       ������������������������       �        ]            �b@        ������������������������       �                      @        B       c       
             �?V��f_�?�            �h@       C       P       	          033�?�S#א��?M            @]@        D       I                   �b@0,Tg��?             E@       E       H                    �?H%u��?             9@       F       G       	          ����?@�0�!��?             1@       ������������������������       �                     ,@        ������������������������       �                     @        ������������������������       �                      @        J       M       	          ����?��.k���?             1@       K       L                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        N       O                   @d@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        Q       `                    w@`2U0*��?4            �R@       R       _                    �?��pBI�?2            @R@       S       ^                    �?`2U0*��?#             I@       T       ]                   �j@���N8�?             E@        U       Z       	          033@z�G�z�?             $@       V       Y                   �a@      �?              @        W       X                   �V@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        [       \       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@        ������������������������       �                      @        ������������������������       �                     7@        a       b                   0c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        d       �       	          033@H���I�?5            �S@       e       h                   @E@���=A�?2             S@        f       g                     P@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        i       v                   �^@�������?-             Q@        j       m                   i@��2(&�?             6@        k       l                     G@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        n       o                   pl@�IєX�?             1@        ������������������������       �                      @        p       q                    �H@�����H�?             "@        ������������������������       �                     @        r       u                    �J@z�G�z�?             @        s       t                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        w       �                    �M@�I� �?             G@       x       y                   �b@�d�����?             C@        ������������������������       �                     (@        z       {                    �?�n_Y�K�?             :@        ������������������������       �                     @        |                          l@�\��N��?             3@        }       ~                   e@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�q�?	             (@       �       �                   �q@�����H�?             "@        ������������������������       �                     @        �       �                    �I@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �c@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ���@      �?           �z@       �       �                    �K@(�7����?�            Py@       �       �                   �`@��2(&�?�            �q@        �       �                    �?�&!��?             �E@       �       �                    X@r٣����?            �@@        ������������������������       �                     �?        �       �                   @c@     ��?             @@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?$�q-�?             :@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        �       �                    �E@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?,�!�?�            `n@        �       �                   0h@���U�?D            �\@       ������������������������       �        C            �[@        ������������������������       �                     @        �       �                    �?(L���?K             `@        ������������������������       �                     @@        �       �       
             �?z�09JX�?<            @X@        �       �                    �?X�<ݚ�?             ;@       �       �                   `a@�û��|�?             7@       �       �                     H@      �?             2@        �       �                   �p@r�q��?             @       ������������������������       �                     @        �       �                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    i@�q�q�?             (@        ������������������������       �                     @        �       �                   �d@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   c@hA� �?)            �Q@        �       �                    �?H%u��?             9@        ������������������������       �                     @        �       �                   @[@r�q��?             2@        ������������������������       �                     @        ������������������������       �        
             .@        ������������������������       �                    �F@        �       �       
             �?�^����?K            �]@       �       �                    �?�z�G��?&             N@       �       �                   `]@      �?             H@        �       �                    @N@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   p`@��i#[�?             E@       �       �                    [@���Q��?             >@        �       �                    @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                    `@D�n�3�?             3@        ������������������������       �                     @        �       �                    �?�q�q�?	             (@        ������������������������       �                     @        �       �                   `_@      �?              @       �       �                   �^@�q�q�?             @       �       �                    �?�q�q�?             @       �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	          033@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     (@        �       �       	             @�j��b�?%            �M@       �       �                   �s@��ϭ�*�?$             M@       �       �                    �L@�1�`jg�?"            �K@        �       �                   @_@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          `ff�?@��8��?             H@       ������������������������       �                     G@        �       �                    �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  }}}}}}�?AAAAAA�?N����4�?-���2�?7`��c.�?��Ug��?�؉�؉�?�;�;�?l(�����?(������?/�袋.�?F]t�E�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?ZZZZZZ�?�������?�?wwwwww�?����X�?����S��?l(�����?�k(����?      �?      �?      �?      �?�������?�������?              �?      �?                      �?�������?ffffff�?UUUUUU�?�������?              �?      �?                      �?      �?        /�袋.�?F]t�E�?              �?�������?�������?              �?      �?                      �?n�%��ʤ?	��wT��?      �?      �?t�E]t�?F]t�E�?              �?      �?      �?      �?                      �?�a�a�?��y��y�?      �?      �?              �?      �?                      �?�0�Ә?9��g9�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?ـl@6 �?�M�&��?              �?      �?        N��)x9�?Y�Cc�?�꡾?��+��+�?1�0��?�y��y��?���Q��?)\���(�?�������?ZZZZZZ�?              �?      �?                      �?�?�������?�q�q�?�q�q�?      �?                      �?      �?      �?      �?                      �?{�G�z�?���Q��?����?���Ǐ�?{�G�z�?���Q��?�a�a�?��y��y�?�������?�������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?                      �?              �?              �?      �?      �?              �?      �?        Q�Ȟ���?^-n����?��P^Cy�?�P^Cy�?      �?      �?              �?      �?        �������?�������?��.���?t�E]t�?333333�?�������?              �?      �?        �?�?      �?        �q�q�?�q�q�?      �?        �������?�������?      �?      �?              �?      �?              �?        Y�B���?Nozӛ��?Cy�5��?y�5���?      �?        ;�;��?ى�؉��?      �?        �5��P�?y�5���?�$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?              �?      �?      �?�u�< �?�)F�?��.���?t�E]t�?֔5eMY�?S֔5eM�?>���>�?|���?              �?      �?      �?UUUUUU�?�������?              �?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?                      �?�_cV�?��L-�?	�#����?p�}��?      �?                      �?⎸#��?w�qG��?      �?        :*����?W?���?�q�q�?r�q��?��,d!�?8��Moz�?      �?      �?�������?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?              �?      �?      �?      �?                      �?���?_�_�?)\���(�?���Q��?      �?        �������?UUUUUU�?              �?      �?              �?        ���?�����?333333�?ffffff�?      �?      �?�������?UUUUUU�?              �?      �?        �<��<��?�a�a�?�������?333333�?F]t�E�?]t�E�?              �?      �?        l(�����?(������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�N��?��/���?����=�?|a���?A��)A�?�־a�?�m۶m��?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ}��NhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM#hzh)h,K ��h.��R�(KM#��h��B�H         >                    �?TU�`��?F           ��@                                  �`@��6}��?v            �f@                                  �J@,�T�6�?B             Z@                     	             @xL��N�?-            �R@                                  �?��pBI�?,            @R@                                   �D@�����?             5@        ������������������������       �                     �?               	       	             �?P���Q�?             4@       ������������������������       �        	             2@        
                           �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      J@        ������������������������       �                     �?                                   e@������?             >@                                 �s@d}h���?             <@                     	          ����?�LQ�1	�?             7@                      
             �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             1@                                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                  �]@V�K/��?4            �S@        ������������������������       �                      @               =       	          `ff@DX�\��?.            �Q@              .       
             �?     ��?)             P@               !                    �?      �?             >@                       	          `ff�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        "       #                    �E@���|���?             6@        ������������������������       �                      @        $       %       	            �?�z�G��?             4@        ������������������������       �                      @        &       '       	          ����?      �?             (@        ������������������������       �                     @        (       )                    @H@      �?              @        ������������������������       �                     �?        *       -                   @b@؇���X�?             @        +       ,                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        /       :                    �?H�V�e��?             A@       0       7                   �s@�r����?             >@       1       2                    �L@ �q�q�?             8@       ������������������������       �        
             *@        3       6                   �d@�C��2(�?             &@        4       5                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        8       9                    t@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ;       <                   Pc@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ?       �       	          ����?l@���?�           ��@        @       {                    �?���6�?�            �u@        A       P       
             �?����X�?f             d@       B       I                   `Z@P��BNֱ?6            �T@        C       D                    Z@�KM�]�?             3@       ������������������������       �                     ,@        E       H                     P@���Q��?             @       F       G       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        J       K                    �?     ��?(             P@       ������������������������       �                      K@        L       M                   �k@ףp=
�?             $@       ������������������������       �                     @        N       O                   �r@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        Q       p                    �?v��:ө�?0            �S@       R       g                   �_@�ՙ/�?'            �O@        S       b       	          ����?���@M^�?             ?@       T       [                   �i@      �?             6@        U       Z                   `]@z�G�z�?             $@       V       Y                   �_@�����H�?             "@        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        \       a                   �^@      �?             (@       ]       `                    �?ףp=
�?             $@        ^       _                    @F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        c       d                    �?�����H�?             "@        ������������������������       �                     @        e       f                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        h       o                    @N@     ��?             @@       i       j                   �d@ףp=
�?             >@       ������������������������       �                     4@        k       l       	          `ffֿ�z�G��?             $@        ������������������������       �                      @        m       n                    �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        q       r                    @I@������?	             .@        ������������������������       �                     @        s       x                   0a@X�<ݚ�?             "@        t       w                    �?z�G�z�?             @       u       v                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        y       z                     L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        |       �       
             �?
QJ�^�?x            �g@        }       �                    @M@�X����?             F@       ~              
             �?�P�*�?             ?@        ������������������������       �                     @        �       �                    �?X�Cc�?             <@        �       �                    �?�z�G��?             $@       �       �                   Pm@�<ݚ�?             "@        �       �                   �i@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          pff�?r�q��?             2@       �       �                    �?      �?             0@       �       �                    �?$�q-�?	             *@        �       �                   �_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?$�q-�?	             *@       ������������������������       �                     "@        �       �                   `c@      �?             @        ������������������������       �                      @        �       �                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �t@ ��֛�?\            @b@       �       �                    �? �}�$>�?Z            �a@        �       �                   0`@�8��8��?	             (@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �       	            �?��"pK�?Q            ``@       ������������������������       �        K             ^@        �       �                    �M@�C��2(�?             &@       �       �                    �?z�G�z�?             @        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?     8�?�             x@        �       �                   �k@V��z4�?K             _@       �       �                    @J@t�7��?'             O@        ������������������������       �        	             ,@        �       �       
             �?�q�q��?             H@        �       �                   �\@      �?              @        ������������������������       �                      @        �       �                   �[@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?R���Q�?             D@       �       �       	          `ff@@4և���?             <@       ������������������������       �                     8@        �       �                    �N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    U@�q�q�?             (@        ������������������������       �                     @        �       �                   �a@      �?              @        �       �                    @L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?V{q֛w�?$             O@       �       �                    @L@:ɨ��?            �@@        �       �                    �?      �?
             0@        ������������������������       �                     @        �       �                   �^@z�G�z�?             $@        ������������������������       �                     �?        �       �       	          ����?�����H�?             "@       �       �                    @H@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�t����?
             1@       �       �                    �?$�q-�?             *@       ������������������������       �                     "@        �       �                   @q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?      �?             @        ������������������������       �                      @        �       �                   Xw@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@�f7�z�?             =@        �       �                    �N@"pc�
�?             &@       ������������������������       �                      @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @r�q��?             2@       ������������������������       �                     &@        �       �                   �a@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �                           @ ����?�            @p@       �       �                   `_@��O���?�            �o@       �       �       
             �?�c!�^�?\            @b@        �       �                   �c@d}h���?             ,@       ������������������������       �        
             $@        �       �                   �X@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   ``@Pa�	�?P            �`@        �       �                    `@���}<S�?              G@       �       �                    _@ >�֕�?            �A@       �       �                   @\@@4և���?             <@        �       �                   �[@�<ݚ�?	             "@       �       �                    Y@      �?              @        �       �                     P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             3@        ������������������������       �                     @        �       �                    �?"pc�
�?	             &@       ������������������������       �                     @        �       �                   �Y@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        0            �U@        �                          �?����?I            @[@       �                         `@0w-!��?C             Y@                                  �?����X�?	             ,@                                0j@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                 �M@���W���?:            �U@                                �?؇���X�?*            �O@                                @M@�3Ea�$�?             G@                   
             �?������?            �B@        	      
                   U@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?�FVQ&�?            �@@                    	          ���@�q�q�?             @        ������������������������       �                     @                                0m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@                    	          ���@X�<ݚ�?             "@                               @_@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     7@                    
             �?X�<ݚ�?             "@                   
             �?����X�?             @        ������������������������       �                      @                                 �L@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        !      "                  �a@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KM#KK��hb�B0  ��Fc*�?y�\���?�!XG��?;ڼOq��?ى�؉��?;�;��?>�S��?L�Ϻ��?���Ǐ�?����?=��<���?�a�a�?              �?ffffff�?�������?      �?              �?      �?      �?                      �?      �?                      �?wwwwww�?�?I�$I�$�?۶m۶m�?��Moz��?Y�B��?      �?      �?              �?      �?              �?        �������?333333�?      �?                      �?              �?�ґ=�?�Z܄��?              �?�]�����?�D+l$�?      �?      �?      �?      �?      �?      �?      �?                      �?F]t�E�?]t�E]�?      �?        333333�?ffffff�?              �?      �?      �?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?iiiiii�?ZZZZZZ�?�������?�?�������?UUUUUU�?      �?        ]t�E�?F]t�E�?�������?�������?              �?      �?              �?              �?      �?              �?      �?              �?      �?              �?      �?                      �?	�2Rl�?y����I�?(��ҁ�?ƯQpZ��?�$I�$I�?�m۶m��?���ˊ��?��FS���?(�����?�k(���?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?     ��?              �?�������?�������?              �?      �?      �?      �?                      �?B�A��?}˷|˷�?�<��<��?�a�a�?�c�1��?�s�9��?      �?      �?�������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�������?�������?      �?        ffffff�?333333�?              �?      �?      �?              �?      �?                      �?�?wwwwww�?              �?�q�q�?r�q��?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?�~�-q�?�c�H;�?]t�E]�?�E]t��?�Zk����?�RJ)���?      �?        �m۶m��?%I�$I��?ffffff�?333333�?9��8���?�q�q�?      �?      �?      �?                      �?      �?                      �?UUUUUU�?�������?      �?      �?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?              �?      �?        ;�;��?�؉�؉�?              �?      �?      �?              �?      �?      �?              �?      �?        {��իW�?�P�B�
�?z��3m��?��^���?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        {k�4w��?qBJ�eD?      �?        ]t�E�?F]t�E�?�������?�������?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?     ��?�s�9��?2�c�1�?��Zk���?SJ)��R�?              �?UUUUUU�?�������?      �?      �?              �?�������?UUUUUU�?              �?      �?        333333�?333333�?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?�������?�������?      �?                      �?      �?        �{����?B!��?e�M6�d�?N6�d�M�?      �?      �?              �?�������?�������?              �?�q�q�?�q�q�?�������?UUUUUU�?              �?      �?              �?        �?<<<<<<�?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?      �?              �?      �?        O#,�4��?a���{�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?        �����?�ȍ�ȍ�?�?�������?Ĉ#F��?t�Ν;w�?۶m۶m�?I�$I�$�?              �?      �?      �?              �?      �?        |���?|���?d!Y�B�?ӛ���7�?�A�A�?��+��+�?�$I�$I�?n۶m۶�?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?              �?F]t�E�?/�袋.�?              �?      �?      �?              �?      �?                      �?j?Y���?&�i?Y�?�p=
ף�?ףp=
��?�$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?      �?                      �?              �?���)kʺ?*kʚ���?�$I�$I�?۶m۶m�?��,d!�?����7��?к����?��g�`��?      �?      �?      �?                      �?|���?>����?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?r�q��?�q�q�?�������?UUUUUU�?              �?      �?                      �?              �?              �?�q�q�?r�q��?�$I�$I�?�m۶m��?              �?�������?333333�?              �?      �?              �?        �������?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJl��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK兔h��B@9         �       
             �?XaG�h�?S           ��@              !                    �?D|U��@�?`           ��@                                   �?v�2t5�?7            �T@                                  b@�+e�X�?"             I@                                  @M@���Q��?             >@                                  i@ҳ�wY;�?             1@        ������������������������       �                     @               	                   �k@      �?
             (@        ������������������������       �                     @        
                          �]@      �?              @        ������������������������       �                     �?                                  �a@؇���X�?             @                                  �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   ]@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     4@                                  �g@     ��?             @@                                   �G@      �?              @        ������������������������       �                     @        ������������������������       �                     @                                  0n@�q�q�?             8@        ������������������������       �                     (@                                   b@�q�q�?	             (@        ������������������������       �                     @                                  �`@      �?              @        ������������������������       �                     @                                    o@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        "       +       	          ����?��)jO�?)           `|@        #       $                   ``@@��!�Q�??            @Z@       ������������������������       �        /             T@        %       &                     D@`2U0*��?             9@        ������������������������       �                     *@        '       *                    j@�8��8��?
             (@        (       )                   �`@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ,       _                    �?
���?�            �u@       -       >                    �?���/��?�            `p@        .       ;                    �?L紂P�?#            �I@       /       2       
             �?�S����?             C@        0       1                   �l@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        3       8                   xr@<���D�?            �@@       4       7       	          ����?XB���?             =@        5       6                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ;@        9       :                   @`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        <       =       	          033�?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ?       @       	          hff�?h+�"��?�            `j@        ������������������������       �                      @        A       T       	          033@ Os���?�             j@       B       E                    \@����� �?o            �e@        C       D                    �?$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        F       S                    �?Уp=
ע?f             d@       G       L                   �e@������?H             \@        H       I       	          033�?��S�ۿ?             >@       ������������������������       �                     .@        J       K                   @e@�r����?	             .@       ������������������������       �                     *@        ������������������������       �                      @        M       R                    �?����ȫ�?4            �T@       N       O                   @a@����e��?)            �P@        ������������������������       �                     @@        P       Q                   �b@г�wY;�?             A@       ������������������������       �                    �@@        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     H@        U       \                   0b@�X�<ݺ?             B@       V       [                    �J@      �?             @@        W       X                   �^@z�G�z�?             @        ������������������������       �                      @        Y       Z                    �I@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        ]       ^       	          `ff@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        `       i                   0`@J�8���?@            �U@        a       h                   P`@�C��2(�?            �@@        b       c                   `d@d}h���?             ,@       ������������������������       �                     $@        d       e                    �?      �?             @        ������������������������       �                     �?        f       g                   �p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        j       {       	          `ff�?      �?*             K@       k       r                    @K@�Gi����?            �B@        l       q       	          ����?�t����?             1@       m       p                   �m@"pc�
�?	             &@        n       o                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        s       v                    �?��Q��?             4@       t       u                   @b@r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        w       x                   �[@      �?              @        ������������������������       �                     @        y       z                   �a@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        |       }                   �b@�t����?             1@        ������������������������       �                     @        ~       �                    �?�eP*L��?
             &@               �                   �k@z�G�z�?             @        �       �                     G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pe@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    I@�>��-��?�            �w@        �       �                   �]@������?             A@        �       �                   �[@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?PN��T'�?             ;@       �       �       	             п�����H�?             2@        ������������������������       �                     �?        �       �                     P@�IєX�?             1@       ������������������������       �        	             ,@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �K@�<ݚ�?             "@        ������������������������       �                     @        �       �                   pa@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?��z��?�            �u@        �       �                    �?䯦s#�?@            �Z@       �       �                    �I@���R�?1            @T@       �       �                    �?�LQ�1	�?             G@        ������������������������       �                     (@        �       �                    �?@�0�!��?             A@        �       �                    @F@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   �d@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   l@`2U0*��?             9@        �       �                   �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             3@        �       �                    �?�xGZ���?            �A@       �       �                    @J@      �?             @@        �       �       	          ����?؇���X�?             @        ������������������������       �                     @        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �L@���Q��?             9@        ������������������������       �                     "@        �       �                   �b@      �?
             0@       �       �                    �O@      �?              @       ������������������������       �                     @        �       �                   `a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @d@ �o_��?             9@       �       �       	          ����?��<b���?             7@        �       �                   n@����X�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             0@        ������������������������       �                      @        �       �                    �?𯁷��?�            @n@        �       �                    �?f1r��g�?            �J@        �       �                    �?�IєX�?             1@        �       �                   �b@r�q��?             @        ������������������������       �                     @        �       �                   �r@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                   �`@tk~X��?             B@        �       �       	          ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    c@��a�n`�?             ?@       ������������������������       �                     9@        �       �                   0c@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @��e�_�?|            �g@       �       �                   @[@�����?r            �e@        �       �                   �b@      �?              @        ������������������������       �                     @        �       �                    c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        k            �d@        �       �                    �?      �?
             0@        ������������������������       �                     "@        �       �                   pg@և���X�?             @        ������������������������       �                     �?        �       �                   �c@�q�q�?             @       �       �                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �A^%���?�Pm4��?�rv��?Xc"=P9�?�ڕ�]��?��+Q��?���Q��?R���Q�?�������?333333�?�������?�������?      �?              �?      �?              �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        ;�;��?�؉�؉�?      �?                      �?              �?      �?      �?      �?      �?      �?                      �?UUUUUU�?�������?      �?        �������?�������?              �?      �?      �?      �?              �?      �?              �?      �?        7%�!6�?Y[�;���?8�8��? �����?              �?{�G�z�?���Q��?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?                      �?              �?A�`���?0�甹��?J�eDP�?���*�?�������?�������?^Cy�5�?(������?�������?333333�?              �?      �?        |���?|���?�{a���?GX�i���?      �?      �?      �?                      �?              �?      �?      �?              �?      �?        ;�;��?�؉�؉�?      �?                      �?H��i�?�� g��?      �?        �$B�e�?����?���"��?����B�?;�;��?�؉�؉�?              �?      �?        333333�?ffffff�?۶m۶m�?I�$I�$�?�?�������?              �?�?�������?              �?      �?        ������?������?|���?�>����?              �?�?�?              �?      �?                      �?              �?�q�q�?��8��8�?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?|a���?�rO#,��?F]t�E�?]t�E�?۶m۶m�?I�$I�$�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?o0E>��?#�u�)��?<<<<<<�?�?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ffffff�?�������?UUUUUU�?�������?      �?                      �?      �?      �?      �?        �������?333333�?              �?      �?        �������?�������?              �?]t�E�?t�E]t�?�������?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�.c��a�?[Ds֠x�?�?xxxxxx�?�$I�$I�?۶m۶m�?              �?      �?        h/�����?&���^B�?�q�q�?�q�q�?      �?        �?�?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?9��8���?              �?�������?333333�?              �?      �?        �2)^ �?v�7[�~�?�����?�V�9�&�?�)O�?��ӭ�a�?��Moz��?Y�B��?      �?        ZZZZZZ�?�������?�q�q�?r�q��?              �?�������?�������?              �?      �?        ���Q��?{�G�z�?�������?UUUUUU�?      �?                      �?      �?        �_�_�?�A�A�?      �?      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?      �?              �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �Q����?
ףp=
�?��Moz��?��,d!�?�m۶m��?�$I�$I�?      �?              �?      �?              �?      �?                      �?      �?        �
�G�?j�V���?�!5�x+�?�x+�R�?�?�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        r�q��?9��8���?�������?�������?              �?      �?        �s�9��?�c�1Ƹ?      �?              �?      �?      �?                      �?t���G'�?p����?&>��?���"�w?      �?      �?      �?              �?      �?              �?      �?              �?              �?      �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ1�)hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKh��B�;         �       
             �?~jÚʞ�?G           ��@              M                    �?���8V�?H           @�@              J                   {@�n���?�            �v@              G                    `R@�dNl`ܾ?�            Pv@                                  �?�1e�3��?�             v@                                   �?z�G�z�?            �F@                                 �e@���!pc�?            �@@        ������������������������       �                     @        	                            K@��X��?             <@        
                           �C@���!pc�?             &@        ������������������������       �                     �?                                  @[@z�G�z�?             $@        ������������������������       �                     �?                                  �q@�����H�?             "@       ������������������������       �                     @                                  �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   i@�IєX�?
             1@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     (@               @                   �b@�]��?�            Ps@                                 �U@�X�
�?�            @r@        ������������������������       �                      @               ?                   `@�=x�?�             r@              "                    �D@��s��?z            �g@               !                    �?      �?             @                                  �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        #       >       	          ����?�g�y��?w            @g@       $       ;                   `_@0G���ջ?E             Z@       %       0                    @O@�nkK�?>             W@       &       /                    �K@ ��PUp�?0            �Q@        '       .                    �?(;L]n�?             >@       (       )                   0l@���7�?             6@       ������������������������       �        
             ,@        *       -       	             �?      �?              @        +       ,                   @`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �D@        1       2                    _@؇���X�?             5@        ������������������������       �                     "@        3       8                   0o@      �?	             (@       4       5                    ]@      �?              @       ������������������������       �                     @        6       7                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        9       :                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        <       =                     L@r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �        2            �T@        ������������������������       �        9             Y@        A       B                    c@�t����?             1@        ������������������������       �                     �?        C       D                     M@      �?             0@       ������������������������       �        	             ,@        E       F                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        H       I                   p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        K       L       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        N       [                    �F@�Q����?h             d@        O       T                   �`@д>��C�?             =@        P       Q                   @`@�q�q�?             @        ������������������������       �                     �?        R       S                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        U       Z                    @ȵHPS!�?             :@       V       Y                   �[@ �q�q�?             8@        W       X                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                      @        \       �       	          `ff�?zVC��?V            ``@       ]       �                    �?�Y �K�?B            @X@       ^       g                    @K@|��?���?(             K@        _       f                   �c@�E��ӭ�?             2@       `       a                   �X@     ��?             0@        ������������������������       �                      @        b       e                   �\@@4և���?	             ,@        c       d                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        h       y                    �?�q�q�?             B@       i       l       	          ����?� �	��?             9@        j       k                   �_@�z�G��?	             $@        ������������������������       �                     @        ������������������������       �                     @        m       n                    �K@������?
             .@        ������������������������       �                      @        o       x                     P@8�Z$���?	             *@       p       q                    �L@����X�?             @        ������������������������       �                      @        r       s       	          ����?���Q��?             @        ������������������������       �                      @        t       u                     N@�q�q�?             @        ������������������������       �                     �?        v       w                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        z       {                    @�C��2(�?	             &@       ������������������������       �                     @        |       �                    �?z�G�z�?             @       }       ~                   @]@�q�q�?             @        ������������������������       �                     �?               �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �[@�ʈD��?            �E@        ������������������������       �                      @        �       �                   `c@������?            �D@       �       �                    �M@�(\����?             D@        �       �                   P`@�IєX�?             1@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     7@        ������������������������       �                     �?        �       �                    �?l��\��?             A@        ������������������������       �                      @        �       �                   �c@      �?             @@       ������������������������       �                     ;@        �       �                   �_@z�G�z�?             @        ������������������������       �                      @        �       �                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?8T���+�?�            �x@       �       �                   @E@̯e<6�?�            0s@        �       �                   �Y@      �?             8@        ������������������������       �                     @        �       �                    �?�t����?             1@       �       �                   �]@$�q-�?             *@       ������������������������       �                      @        �       �       	             пz�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@�����Z�?�            �q@        �       �                   Hp@@���?-�?X            �a@       ������������������������       �        A            �Z@        �       �                    @�8��8��?             B@       �       �                   xp@г�wY;�?             A@        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                      @        �       �                    �L@`	�<��?\            �a@       �       �                   �l@_k,D	�?P            �]@        �       �                   �e@@3����?%             K@       ������������������������       �                     D@        �       �                    �?@4և���?             ,@        �       �                   0f@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             $@        �       �                   �f@      �?+             P@       �       �                    �?�����H�?*            �O@        �       �                    `@X�Cc�?	             ,@        �       �                   �c@r�q��?             @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   0c@@9G��?!            �H@        ������������������������       �                     �?        �       �                    �?@��8��?              H@        �       �                    �K@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     C@        ������������������������       �                     �?        �       �                   �r@\X��t�?             7@       �       �                    �?      �?             0@        �       �                    \@      �?              @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �c@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?և���X�?=            �V@        �       �                   �Z@ףp=
�?             >@        ������������������������       �                      @        �       �                   `T@h�����?             <@        ������������������������       �                     �?        ������������������������       �                     ;@        �       �                   �]@Nd^����?*            �N@        ������������������������       �        
             ,@        �       �                    �?JJ����?             �G@       �       �                     P@��<b���?             7@       �       �                    �J@�KM�]�?             3@        ������������������������       �                      @        �       �                    �K@"pc�
�?             &@        ������������������������       �                     �?        �       �                    �M@ףp=
�?             $@        �       �                    @M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	             @r�q��?             8@       �       �                    U@�LQ�1	�?             7@        ������������������������       �                     �?        �       �       	          ����?�C��2(�?             6@        �       �                   �d@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             1@        ������������������������       �                     �?        �t�b�<     h�h)h,K ��h.��R�(KK�KK��hb�B�  g�����?L��/��?�J��J��?K��J���?r�qǱ?r�q��?5~5~�?^9�]9��?W'u_�?�/���?�������?�������?t�E]t�?F]t�E�?              �?%I�$I��?n۶m۶�?F]t�E�?t�E]t�?              �?�������?�������?              �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?�?�?      �?      �?      �?                      �?              �?              �?��,�?p�14���?�1bĈ�?w�ܹs��?      �?        ����?�?8���?�X�0Ҏ�?q�����?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�B!��?��{���?�؉�؉�?vb'vb'�?d!Y�B�?�Mozӛ�?��V،?��ۥ���?�?�������?F]t�E�?�.�袋�?              �?      �?      �?      �?      �?              �?      �?                      �?              �?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?                      �?              �?�?<<<<<<�?      �?              �?      �?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?a���{�?|a���?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ��N��N�?�؉�؉�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?V���g�?ձ�6Ls�?����?���
|q�?{	�%���?	�%����?�q�q�?r�q��?      �?      �?              �?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?�������?�������?�Q����?)\���(�?333333�?ffffff�?      �?                      �?wwwwww�?�?              �?;�;��?;�;��?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        F]t�E�?]t�E�?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?�}A_з?A_���?      �?        ������?p>�cp�?�������?333333�?�?�?      �?      �?              �?      �?                      �?              �?      �?        �������?------�?      �?              �?      �?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�~r!�?���6z�?���t�?�j�Z�?      �?      �?              �?�������?�������?�؉�؉�?;�;��?      �?        �������?�������?      �?                      �?              �?��*��?�Co߫�?^����R�?H���@��?      �?        UUUUUU�?UUUUUU�?�?�?              �?      �?                      �?o����?E�)͋?�?����/��?��c+���?���Kh�?h/�����?      �?        n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?              �?      �?�q�q�?�q�q�?%I�$I��?�m۶m��?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        ������?9/���?              �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?                      �?!Y�B�?��Moz��?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?�$I�$I�?۶m۶m�?�������?�������?              �?�m۶m��?�$I�$I�?              �?      �?        ���:�?�u�y���?              �?��
br�?x6�;��?��Moz��?��,d!�?(�����?�k(���?              �?F]t�E�?/�袋.�?      �?        �������?�������?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?�������?UUUUUU�?��Moz��?Y�B��?              �?]t�E�?F]t�E�?333333�?�������?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�u�ThG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM#hzh)h,K ��h.��R�(KM#��h��B�H         2                    _@X�<ݚ�?8           ��@                                   �?$�{�F"�?j             e@                                  �?�C��2(�?K            @^@                                   �?H.�!���?              I@              
       	             �?�חF�P�?             ?@                                  �`@@4և���?
             ,@       ������������������������       �                     &@               	                   pb@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  `@������?             1@       ������������������������       �        	             (@                      	             @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                                  @]@�����?	             3@                                   �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @                      
             �?8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �        +            �Q@               #       
             �?�q�q�?             H@                      	             @��S�ۿ?             >@                                  @O@h�����?             <@       ������������������������       �        
             1@                                   �O@�C��2(�?             &@                                  �\@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        !       "                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        $       +                    �?�q�q�?             2@       %       &                    ^@      �?              @        ������������������������       �                     @        '       (                   @_@      �?             @        ������������������������       �                      @        )       *                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                     M@�z�G��?             $@        ������������������������       �                      @        .       1       	             �?      �?              @       /       0                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        3       �                    �?������?�           h�@       4                           @L@��$�ƹ�?"           @}@       5       J                    �?@�0�!��?�            0t@        6       =       
             �?yÏP�?3            �T@        7       <                   �e@6YE�t�?            �@@       8       9       	          ����?��S�ۿ?             >@       ������������������������       �                     2@        :       ;                    �?r�q��?	             (@        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        >       I                    �G@؇���X�?            �H@       ?       H                   @_@ �o_��?             9@        @       A                   �i@�q�q�?	             (@        ������������������������       �                     @        B       C                    �?X�<ݚ�?             "@        ������������������������       �                     �?        D       E                   �a@      �?              @        ������������������������       �                     @        F       G                    �E@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        ������������������������       �                     8@        K       h       	          ����?��w]j<�?�             n@       L       ]       
             �?����!p�?w             f@        M       V                   pd@���Q��?             4@        N       O                    �?�q�q�?             "@        ������������������������       �                     �?        P       U                    @      �?              @       Q       R                    �B@�q�q�?             @        ������������������������       �                      @        S       T                    @G@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        W       \                    �?"pc�
�?             &@       X       Y                    �?ףp=
�?             $@        ������������������������       �                     @        Z       [                   �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ^       g                    �?�(�Tw�?g            �c@       _       `                   @n@ ��ʻ��?X             a@       ������������������������       �        5            @T@        a       f                   0c@h㱪��?#            �K@        b       c                    �?�t����?             1@        ������������������������       �                     @        d       e                   �n@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     C@        ������������������������       �                     4@        i       p                    �?�����D�?!            @P@        j       o       	          ����?h�����?             <@        k       l       	          pff�?r�q��?             @        ������������������������       �                     @        m       n                    �F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             6@        q       r                   Pa@V������?            �B@        ������������������������       �                     $@        s       v                   @m@�5��?             ;@        t       u                     G@      �?              @        ������������������������       �                      @        ������������������������       �                     @        w       z       	          ����?�d�����?             3@        x       y                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        {       |                    @�C��2(�?             &@       ������������������������       �                     "@        }       ~                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?20J�Ws�?W             b@        �       �                    �?�G�5��?(            @Q@       �       �                   Xv@j�q����?             I@       �       �       
             �?�LQ�1	�?             G@       ������������������������       �                     ?@        �       �                   �b@���Q��?	             .@        ������������������������       �                     @        �       �                    �L@ףp=
�?             $@        �       �                   0d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @O@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �N@D�n�3�?             3@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �b@���|���?
             &@        �       �                    @���Q��?             @       �       �                   P`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @r�q��?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �h@\�Uo��?/             S@        �       �                    �?�����H�?             2@        ������������������������       �                      @        �       �                   �`@z�G�z�?             $@        ������������������������       �                     �?        �       �                   �`@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   q@l��[B��?#             M@       �       �                    �?�K��&�?            �E@        �       �                    @z�G�z�?             @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Hp@p�ݯ��?             C@       �       �                   `k@l��[B��?             =@        �       �       
             �?�����H�?             "@       ������������������������       �                     @        �       �                    j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �k@��Q��?             4@        ������������������������       �                     @        �       �                   0o@��
ц��?	             *@       �       �                   �`@�<ݚ�?             "@        ������������������������       �                     @        �       �                    @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?z�G�z�?	             .@       ������������������������       �                     $@        �       �                    Z@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �                         �b@hX͇���?�            �q@       �       �                    �?6C�d�?�            �o@        �       �                   �g@���"͏�?            �B@        ������������������������       �                      @        �       �       
             �?z�G�z�?            �A@       �       �                   hu@6YE�t�?            �@@       �       �                   @m@ףp=
�?             >@        �       �                    �?      �?              @       �       �       	             �?      �?             @        ������������������������       �                     �?        �       �                   `a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     6@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �                         Hq@�g��?�            �j@       �                          @n�3���?Z             c@       �       �       	          ����?v���a�?W            @b@        �       �                    �?r�qG�?             H@        �       �       
             �?�t����?
             1@       ������������������������       �                     ,@        �       �                    o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �o@�g�y��?             ?@       �       �                   �\@�q�q�?             5@        ������������������������       �                     @        �       �                   `Z@�<ݚ�?             2@        �       �                    �?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             &@        �       �                    �?z�G�z�?             $@       �       �                    �?�����H�?             "@       �       �                    Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?ؗp�'ʸ?:            �X@        �       �                   �Z@�t����?
             1@        ������������������������       �                     �?        �       �       
             �?      �?	             0@       �       �                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �J@ 7���B�?0            @T@        �       �                   �_@؇���X�?
             ,@        �       �                   �^@�q�q�?             @        ������������������������       �                     @        �       �                   @]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �                         �\@�\=lf�?&            �P@        �                            N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        $            @P@                                �j@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                �\@�i�y�?(            �O@                                 �R@�t����?             1@                                �?      �?             0@       	            	             �?$�q-�?             *@        
                        �s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             &@        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     G@                                 `@П[;U��?             =@                    
             �?�q�q�?
             .@                                �?�eP*L��?             &@        ������������������������       �                      @                                 @C@�q�q�?             "@        ������������������������       �                     @                                @c@      �?             @        ������������������������       �                      @                                 �F@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              "                  0p@d}h���?             ,@             !                   �?�z�G��?	             $@                                  M@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM#KK��hb�B0  �q�q�?r�q��?��WV��?�	j*D�?F]t�E�?]t�E�?)\���(�?�(\����?��RJ)��?�Zk����?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?      �?                      �?�?xxxxxx�?              �?�������?�������?      �?                      �?^Cy�5�?Q^Cy��?UUUUUU�?UUUUUU�?      �?                      �?;�;��?;�;��?              �?      �?                      �?�������?�������?�?�������?�$I�$I�?�m۶m��?              �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?      �?      �?                      �?ffffff�?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        -ьt�\�?�]�F�?��~��~�?#0#0�?ZZZZZZ�?�������?W�v%jW�?Q��+Q�?e�M6�d�?'�l��&�?�?�������?              �?UUUUUU�?�������?      �?                      �?      �?        ۶m۶m�?�$I�$I�?
ףp=
�?�Q����?�������?�������?              �?r�q��?�q�q�?      �?              �?      �?      �?        �������?�������?      �?                      �?      �?              �?        �.�.�?�^�^�?/�袋.�?]t�E�?333333�?�������?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?/�袋.�?F]t�E�?�������?�������?      �?        �������?UUUUUU�?      �?                      �?              �?p��o���?�A�A�?�������?�?      �?        ־a���?��)A��?<<<<<<�?�?      �?        /�袋.�?F]t�E�?              �?      �?              �?              �?        z�z��?z�z��?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �g�`�|�?o0E>��?      �?        h/�����?/�����?      �?      �?      �?                      �?Cy�5��?y�5���?      �?      �?              �?      �?        ]t�E�?F]t�E�?      �?              �?      �?              �?      �?        �Ő��?z�!���?�%~F��?��v`��?
ףp=
�?=
ףp=�?Y�B��?��Moz��?              �?�������?333333�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?(������?l(�����?      �?      �?              �?      �?        ]t�E]�?F]t�E�?�������?333333�?      �?      �?      �?                      �?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?�5��P^�?6��P^C�?�q�q�?�q�q�?      �?        �������?�������?              �?�q�q�?�q�q�?              �?      �?        ���=��?GX�i���?���)k��?��)kʚ�?�������?�������?      �?      �?      �?                      �?      �?        Cy�5��?^Cy�5�?GX�i���?���=��?�q�q�?�q�q�?              �?      �?      �?              �?      �?        �������?ffffff�?      �?        �؉�؉�?�;�;�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�������?      �?        �������?333333�?      �?                      �?��\���?��h����?�4M�4M�?˲,˲,�?*�Y7�"�?v�)�Y7�?      �?        �������?�������?e�M6�d�?'�l��&�?�������?�������?      �?      �?      �?      �?              �?333333�?�������?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �=��C�?��U��?�k(����?�5��P�?�4iҤI�?ٲe˖-�?�������?�������?�?<<<<<<�?              �?UUUUUU�?UUUUUU�?      �?                      �?��{���?�B!��?UUUUUU�?UUUUUU�?      �?        �q�q�?9��8���?�$I�$I�?۶m۶m�?              �?      �?                      �?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?              �?                      �?����X�?�S�r
^�?�?<<<<<<�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?h/�����?	�%����?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?g��1��?"=P9���?      �?      �?      �?                      �?              �?�������?UUUUUU�?      �?                      �?AA�?�������?�?<<<<<<�?      �?      �?;�;��?�؉�؉�?      �?      �?      �?                      �?              �?              �?      �?                      �?�{a���?��=���?UUUUUU�?UUUUUU�?]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?                      �?              �?I�$I�$�?۶m۶m�?ffffff�?333333�?9��8���?�q�q�?      �?                      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ݂#yhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@>         .                    �?��.k���?E           ��@                      
             �?�y���?~            �h@                                  �Q@V�K/��?3            �S@        ������������������������       �                     &@                                  �a@h+�v:�?-             Q@                                  �?R�}e�.�?!             J@                                  �?�û��|�?             7@                                  �?�\��N��?             3@        	       
                   �`@؇���X�?             @       ������������������������       �                     @                      	          033@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  �g@      �?
             (@        ������������������������       �                     �?                                   �?"pc�
�?	             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     =@                      	          ����?      �?             0@        ������������������������       �                     @                                   @H@$�q-�?
             *@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@               !                    T@P���Q�?K             ^@                                   @b@      �?             @                                 �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        "       )                    �?P�Lt�<�?H            �\@       #       (                    �?�����??            @Y@        $       %                   �b@P���Q�?             4@       ������������������������       �        
             1@        &       '                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        3            @T@        *       +                     L@8�Z$���?	             *@        ������������������������       �                     @        ,       -                    �M@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        /       �                    �?�ه�F�?�           x�@       0       c       
             �?�N_��?�            px@        1       `                    f@x��}�?f            �d@       2       E                    �?X�If%��?]            �b@       3       6                   �Q@P��BNֱ?4            �T@        4       5       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        7       @                   �r@F|/ߨ�?2            @T@       8       9       	          ����?�"w����?.             S@       ������������������������       �                     D@        :       ?                    �M@������?             B@        ;       <                   �`@$�q-�?	             *@       ������������������������       �                      @        =       >                    @M@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     7@        A       B       	          ����?z�G�z�?             @        ������������������������       �                     @        C       D                     O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        F       _                   Pq@�4��?)            @P@       G       R                    �?l`N���?#            �J@        H       Q                   �c@p�ݯ��?             3@       I       L                   0c@��
ц��?	             *@       J       K                     M@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        M       N                   �c@����X�?             @        ������������������������       �                     @        O       P                   �k@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        S       V                    �?�t����?             A@        T       U                   o@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        W       X       	             �?���}<S�?             7@       ������������������������       �        	             0@        Y       ^                   `c@����X�?             @       Z       [                   0b@r�q��?             @        ������������������������       �                     @        \       ]                   Pb@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        a       b                   `e@@�0�!��?	             1@        ������������������������       �                     @        ������������������������       �                     ,@        d       y                    �?D+ҭb��?�            @l@        e       x                    �?#z�i��?            �D@       f       g                     D@`՟�G��?             ?@        ������������������������       �                     @        h       i                   @\@|��?���?             ;@        ������������������������       �                     @        j       k                   `\@�q�q�?             5@        ������������������������       �                     @        l       w                   Pq@      �?             ,@       m       v                     M@���|���?
             &@       n       u       	          833�?      �?              @       o       p                   �m@և���X�?             @        ������������������������       �                     @        q       r                    �F@      �?             @        ������������������������       �                      @        s       t       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        z       �                    �?T}_���?v             g@       {       �                   @[@D���D|�?e            �c@        |                          @c@���Q��?             @        }       ~                    �G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    _@xJ��b,�?a            @c@        ������������������������       �                    �H@        �       �                    �?�#-���?B            @Z@       �       �                   �_@ܷ��?��?9            �U@        �       �                    �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @��(\���?5             T@       �       �                    @N@�kb97�?3            @S@       �       �                   �b@��?^�k�?.            �Q@       ������������������������       �        (            �N@        �       �                   `n@�<ݚ�?             "@       �       �                   @k@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �c@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                     O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             2@        �       �                    �?��
ц��?             :@       �       �                   @^@X�<ݚ�?             2@        ������������������������       �                     @        �       �                   �O@�q�q�?
             .@        ������������������������       �                     @        ������������������������       �                     $@        �       �                    �?      �?              @       �       �       	          (33�?և���X�?             @       �       �                   �a@      �?             @        ������������������������       �                      @        �       �                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   `d@�p ��?�            �t@       �       �                   P`@�6@�?�            �s@       �       �                   �[@��M�'�?�            �k@        �       �                     E@���7�?2             V@        ������������������������       �                      @        �       �                   �[@ qP��B�?1            �U@        �       �                    �?z�G�z�?             $@        �       �       	          ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        -             S@        �       �       
             �?�\�)G�?\            �`@       �       �       	          ����?�S���?S             ^@       �       �       	          033�?l��\��?/             Q@       �       �                    @M@�nkK�?"             G@       ������������������������       �                     >@        �       �                   p`@      �?             0@        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �E@"pc�
�?             6@        �       �                    b@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             0@       �       �                   �j@      �?              @        �       �                   �]@�q�q�?             @        ������������������������       �                     �?        �       �                   pe@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   8p@ pƵHP�?$             J@       ������������������������       �                     A@        �       �                    @K@�X�<ݺ?             2@        �       �                   �q@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   @b@���Q��?	             .@       �       �                   @]@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   �^@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�q�Q�?<             X@       �       �                   �Z@:�&���?0            �S@        ������������������������       �                     @        �       �                   �m@$G$n��?.            �R@       �       �       
             �?R���Q�?             D@       �       �                   �\@�����H�?             ;@        �       �                   �j@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     3@        �       �                    b@��
ц��?             *@       �       �                   a@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    c@г�wY;�?             A@       ������������������������       �                     ;@        �       �                    q@؇���X�?             @        ������������������������       �                     @        �       �                   �q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    Y@      �?             2@        ������������������������       �                     @        �       �                   m@���Q��?             .@        ������������������������       �                     @        �       �                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �C@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �?�������?�큍��?
H�Ʌ��?�ґ=�?�Z܄��?              �?�������?xxxxxx�?'vb'vb�?�;�;�?��,d!�?8��Moz�?�5��P�?y�5���?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?      �?      �?        F]t�E�?/�袋.�?      �?                      �?              �?      �?              �?      �?      �?        ;�;��?�؉�؉�?      �?      �?              �?      �?                      �?ffffff�?�������?      �?      �?      �?      �?              �?      �?                      �?���k(�?(�����?�tj��?��be�F�?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ;�;��?;�;��?      �?        �m۶m��?�$I�$I�?              �?      �?        =ʸ�D��?�#�]��?:���?���(��?A��)A�?pX���o�?�Y7�"��?�)�Y7��?���ˊ��?��FS���?      �?      �?      �?                      �?�����H�?�Hx�5�?(�����?Cy�5��?              �?�q�q�?�q�q�?;�;��?�؉�؉�?              �?�������?�������?              �?      �?                      �?�������?�������?              �?      �?      �?              �?      �?        �Z��Z��?�R+�R+�?
�[���?�R���?^Cy�5�?Cy�5��?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?F]t�E�?t�E]t�?      �?                      �?d!Y�B�?ӛ���7�?              �?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?ZZZZZZ�?�������?              �?      �?        O-�����?�JO-���?�+Q��?ە�]���?�1�c��?�s�9��?      �?        	�%����?{	�%���?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?]t�E]�?F]t�E�?      �?      �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?              �?      �?      �?                      �?      �?              �?                      �?      �?        Y�����?<��ӿ?*Z8B��?�.=�ﵱ?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ��8+?!�?5�wL�?      �?        �A�A�?_�_�?��=���?a���{�?�$I�$I�?۶m۶m�?              �?      �?        �������?333333�?�Y�	qV�?�cj`?_�_��?�A�A�?      �?        9��8���?�q�q�?333333�?�������?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �;�;�?�؉�؉�?r�q��?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?              �?      �?                      �?      �?        ��+Q��?Q��+Q�?�*u��?^�b;���? �����?|�m��?F]t�E�?�.�袋�?      �?        �}A_З?��}A�?�������?�������?      �?      �?              �?      �?                      �?              �?n�Q�ߦ�?�Ε$��?�����ݭ?""""""�?�������?------�?d!Y�B�?�Mozӛ�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?/�袋.�?      �?      �?              �?      �?              �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?;�;��?'vb'vb�?              �?�q�q�?��8��8�?�q�q�?�q�q�?      �?                      �?              �?�������?333333�?r�q��?�q�q�?      �?        �������?�������?              �?      �?        UUUUUU�?�������?              �?      �?        �������?UUUUUU�?�o��o��?�A�A�?      �?        ���L�?к����?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?                      �?�؉�؉�?�;�;�?      �?      �?      �?                      �?      �?        �?�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?      �?              �?333333�?�������?      �?              �?      �?              �?      �?        �q�q�?�q�q�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�^�@hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK酔h��B@:         �       
             �?X�<ݚ�?>           ��@              ?                    �?�#l��?@           �@              >                   `f@@4և���?�            �v@                                 �U@�IQu`�?�            �v@        ������������������������       �                     �?               /                   Pa@Ȝ�Ѫ2�?�            pv@              .                    �?��H���?|             h@                                 �h@��l�5�?Y            `a@        	       
                    _@�Ń��̧?             E@       ������������������������       �                     8@                                  �_@�X�<ݺ?             2@                                   �P@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@                                  0i@z�09JX�?>            @X@                                  �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?               )                   �b@t/*�?;            �W@              $                    �?�Zl�i��?4            @T@                                 �Z@ >�֕�?-            �Q@                      	              @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                  Xp@�����?*            �P@       ������������������������       �                    �@@               #                    `@l��\��?             A@                                  xp@      �?             (@        ������������������������       �                     �?                                   Pr@"pc�
�?             &@       ������������������������       �                     @        !       "                    @D@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     6@        %       &                   �j@���|���?             &@        ������������������������       �                      @        '       (                   �l@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        *       +                   pd@�n_Y�K�?             *@        ������������������������       �                     @        ,       -       	          @33�?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        #             K@        0       =                    �?��'�`�?_            �d@       1       <                    @H@�T�~~4�?C            @]@        2       ;                   �m@�����?             5@        3       4       	             �?      �?              @        ������������������������       �                      @        5       6                    b@�q�q�?             @        ������������������������       �                      @        7       8                     F@      �?             @        ������������������������       �                     �?        9       :       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �        4             X@        ������������������������       �                    �H@        ������������������������       �                     @        @       �                    �?֭��F?�?c            �a@       A       �                    `Q@��o	��?R             ]@       B       Q                    �?xO�a���?N            @[@        C       P       	          ����?�'�`d�?            �@@       D       I                   `m@p�ݯ��?             3@       E       H       	          ����?"pc�
�?             &@       F       G                    T@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        J       K                    �?      �?              @        ������������������������       �                     @        L       O                   �a@���Q��?             @       M       N                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        R       e                    �?&:~�Q�?9             S@        S       T                   �[@l��[B��?             =@        ������������������������       �                     @        U       d                    �?      �?             8@       V       W                   0g@�\��N��?             3@        ������������������������       �                     @        X       _                    @     ��?             0@        Y       Z       	          833�?      �?              @        ������������������������       �                     �?        [       \                    `@؇���X�?             @       ������������������������       �                     @        ]       ^       	          hff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        `       c                    �?      �?              @       a       b                   pq@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        f                          �f@�7����?$            �G@       g       t                    �?��Hg���?"            �F@        h       o                    �K@�n_Y�K�?             *@       i       n                     G@�<ݚ�?             "@       j       k                   �a@���Q��?             @        ������������������������       �                     �?        l       m                   0m@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        p       s                    �?      �?             @       q       r                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        u       v                   `X@     ��?             @@        ������������������������       �                     �?        w       ~                   �b@�חF�P�?             ?@       x       y                    �?�r����?             >@       ������������������������       �                     .@        z       }       	          ����?������?	             .@       {       |       	             �?X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@        �       �                   @E@���j��?�            �y@        �       �                   �`@^l��[B�?             M@       �       �       	            �?      �?             @@        �       �                    `R@r�q��?             (@       �       �                    �?�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                   �_@      �?             @        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          033�?ףp=
�?	             4@       ������������������������       �                     1@        �       �                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@ ��WV�?             :@       ������������������������       �        	             0@        �       �       	          hff�?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?�Z��L��?�            0v@        �       �       	            �?���3�E�?<             Z@       �       �                   �b@8�Z$���?.            �S@       ������������������������       �                     F@        �       �                    @C@ҳ�wY;�?             A@        ������������������������       �                     "@        �       �                   0c@�q�����?             9@        ������������������������       �                     @        �       �                    �N@8�A�0��?             6@       �       �                    �?      �?             2@        �       �                    b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?և���X�?
             ,@       �       �                   @Z@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                    k@�q�q�?             @        ������������������������       �                      @        �       �                   �_@      �?             @        ������������������������       �                     �?        �       �                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �l@z�G�z�?             @       �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�	j*D�?             :@        ������������������������       �                     @        �       �                    `P@ףp=
�?             4@       ������������������������       �        	             ,@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @0i��?�            `o@       �       �                   0h@��x$�?�            �l@       �       �                   �s@0���U'�?�            @l@       �       �                    �?@�n���?�            �i@        ������������������������       �        1             T@        �       �       	            �? ������?V            �_@       �       �                    �?����r�?I            �[@        �       �                   `b@@4և���?
             ,@       ������������������������       �                     (@        �       �                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        ?             X@        �       �                    @L@      �?             0@       ������������������������       �                      @        �       �                    �M@      �?              @        �       �                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �s@R���Q�?             4@        ������������������������       �                     �?        �       �                    �N@�KM�]�?             3@       ������������������������       �        	             ,@        �       �                   �u@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �D@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    @M@��s����?             5@       ������������������������       �        	             .@        �       �                    ^@�q�q�?             @        ������������������������       �                     �?        �       �       	          ����?z�G�z�?             @        ������������������������       �                     @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �q�q�?r�q��?��be�F�?�I��A��?�$I�$I�?n۶m۶�?��I��I�?�`�`�?      �?        �V�*�?�Z�^� �?�ҡ�3�?��+����??ZMB�?p�l�:��?�a�a�?��<��<�?              �?�q�q�?��8��8�?      �?      �?              �?      �?                      �?W?���?:*����?UUUUUU�?UUUUUU�?      �?                      �?W�+���?�;����?�����H�?�"e����?�A�A�?��+��+�?UUUUUU�?UUUUUU�?              �?      �?        ���@��?g��1��?              �?�������?------�?      �?      �?      �?        F]t�E�?/�袋.�?              �?�������?333333�?              �?      �?                      �?F]t�E�?]t�E]�?      �?        �q�q�?9��8���?              �?      �?        ;�;��?ى�؉��?      �?        UUUUUU�?�������?              �?      �?                      �?��k���?1P�M��?���??�s?�s�?�a�a�?=��<���?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?      �?        br1���?�F}g���?������?���{�?��]8��?��p�?6�d�M6�?'�l��&�?^Cy�5�?Cy�5��?/�袋.�?F]t�E�?�������?�������?              �?      �?                      �?      �?      �?              �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �k(����?�k(���?GX�i���?���=��?      �?              �?      �?�5��P�?y�5���?              �?      �?      �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?      �?۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?G}g����?]AL� &�?��I��I�?؂-؂-�?ى�؉��?;�;��?�q�q�?9��8���?�������?333333�?              �?      �?      �?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?        ��RJ)��?�Zk����?�?�������?              �?�?wwwwww�?�q�q�?r�q��?              �?      �?                      �?      �?              �?        �$I�$I�?۶m۶m�?      �?                      �?              �?�f���i�?kdv�X�?��=���?�=�����?      �?      �?�������?UUUUUU�?9��8���?�q�q�?              �?      �?      �?      �?      �?      �?      �?      �?                      �?      �?              �?              �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?O��N���?              �?�������?�������?      �?                      �?���.�d�?��Vؼ?O��N���?b'vb'v�?;�;��?;�;��?      �?        �������?�������?      �?        �p=
ף�?���Q��?              �?颋.���?/�袋.�?      �?      �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?      �?        ;�;��?vb'vb'�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�/� ���?���e�?�aܯK*�?��s���?-����J�?Vzja���?\mMw��?��,�?      �?        ��}��}�?AA�?�oX����?��)A��?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?              �?              �?      �?      �?              �?      �?      �?      �?      �?                      �?      �?        333333�?333333�?              �?�k(���?(�����?      �?        333333�?�������?              �?      �?              �?      �?      �?                      �?z��y���?�a�a�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?      �?                      �?�t�bub��"     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ,ǁhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK煔h��B�9         "                   �_@�7i���?L           ��@                                   �?,sI�v�?n            �f@                                   �?ڤ���?2            @T@                                   �N@�5��?             ;@                                  @D@�8��8��?
             (@        ������������������������       �                     �?        ������������������������       �        	             &@               	       	          ����?�q�q�?             .@        ������������������������       �                     @        
                          @L@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?                      
             �?r�q��?              K@        ������������������������       �                     @                      
             �?�t����?            �I@                                  �?��Y��]�?            �D@       ������������������������       �                     ?@                                    M@ףp=
�?             $@       ������������������������       �                     @                                   �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  0a@      �?             $@        ������������������������       �                     @                      	             �?r�q��?             @        ������������������������       �                     @                                   �I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?��F�D�?<            �X@       ������������������������       �        ,             R@                !       	             @�>����?             ;@       ������������������������       �                     9@        ������������������������       �                      @        #       �       	          `ff�?⧓Yd��?�           �@       $       ?       
             �?�U���S�?           �y@        %       .                    �?�L�lRT�?E            �V@        &       +                   `a@"pc�
�?             6@       '       *                    @N@�����H�?             2@       (       )                    �?�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �                     �?        ,       -                   �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        /       0       	          ����?H�V�e��?4             Q@       ������������������������       �        "            �E@        1       6                   �a@� �	��?             9@        2       5                   �`@�z�G��?	             $@       3       4                   �p@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        7       8       
             �?������?	             .@        ������������������������       �                     @        9       >                    �?���|���?             &@       :       ;                    �?�<ݚ�?             "@       ������������������������       �                     @        <       =                     J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        @       S                   �]@��[��^�?�            0t@        A       H                   �b@^��4m�?+            �R@       B       G       	          pff�?�X�<ݺ?             B@       C       D                    �?��?^�k�?            �A@       ������������������������       �                    �@@        E       F                   @[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        I       J                    �?�s��:��?             C@        ������������������������       �                     *@        K       R                    �?`�Q��?             9@       L       O                    �?��+7��?             7@        M       N                   �e@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        P       Q                   c@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        T       o                    �?��仞�?�             o@        U       b                    �?��a�n`�?'             O@        V       ]                    �?�G�z��?             4@       W       X                   0n@�eP*L��?             &@        ������������������������       �                     @        Y       \                    d@      �?              @        Z       [       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ^       a                    �?X�<ݚ�?             "@       _       `                   �`@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        c       d                    �?@4և���?             E@        ������������������������       �                     $@        e       l                   �b@     ��?             @@       f       k                   pf@XB���?             =@        g       j                    �?�q�q�?             @       h       i                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        m       n                   po@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        p       �                   �g@��R�x��?{            `g@       q       ~                    @f�1�?z             g@       r       y                    �O@0���ަ?r            �e@       s       t                   �`@�=
ףp�?j             d@       ������������������������       �        E            �Z@        u       x                    a@�O4R���?%            �J@        v       w                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        #            �I@        z       {                    �?z�G�z�?             .@       ������������������������       �                     $@        |       }                    �P@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @               �                   hp@z�G�z�?             $@       �       �                   �k@�����H�?             "@        �       �       	            �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��:"��?�            Pt@       �       �                    �?X�;�^o�?�            �k@        �       �                   ``@����>�?            �B@        �       �                    s@�eP*L��?             &@       �       �                   �q@�q�q�?             "@       �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?8�Z$���?             :@       �       �       	          ����?H%u��?             9@        �       �       	          ����?      �?              @       �       �                    �H@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     �?        �       �                    f@\#r��?s            �f@       �       �                    �? ]�� ��?r            �f@        �       �                   ``@      �?             <@        ������������������������       �                     *@        �       �                    b@��S���?             .@       �       �                    a@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �F@�IєX�?b             c@        �       �       	             @      �?             4@       �       �                     E@�t����?             1@       �       �                    `@      �?              @        �       �                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        �       �                   �\@Pns��ޭ?U            �`@        �       �                   Pk@؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        �       �                    @M@ ����?M            �]@       ������������������������       �        .             R@        �       �                   �b@`�q�0ܴ?            �G@       ������������������������       �                    �F@        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?<W#.m��??            @Z@        �       �                    �?(N:!���?            �A@        ������������������������       �                     $@        �       �                    �H@�J�4�?             9@        �       �                   �b@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?�KM�]�?             3@       �       �                   @q@r�q��?             (@       ������������������������       �                      @        �       �                   @_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �l@���Q��?*            �Q@        �       �                     N@J�8���?             =@       �       �                   �a@��s����?             5@        �       �       	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   f@�����H�?	             2@        ������������������������       �                     �?        �       �                   �k@�IєX�?             1@       ������������������������       �                     (@        �       �       	          ���@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �O@      �?              @        ������������������������       �                     @        �       �                   �j@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �B@��P���?            �D@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @J@4?,R��?             B@        ������������������������       �                     (@        �       �                   hq@�q�q�?             8@       �       �                   @^@�q�q�?	             .@        ������������������������       �                     @        �       �                   �b@�eP*L��?             &@       �       �                    �L@      �?              @        �       �                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  }}}}}}�?AAAAAA�?��I��I�?l�l��?X�<ݚ�?����H�?/�����?h/�����?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?]t�E�?F]t�E�?      �?                      �?UUUUUU�?�������?      �?        �?<<<<<<�?������?8��18�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        [�R�֯�?j�J�Z�?              �?h/�����?�Kh/��?              �?      �?        ��k5c�?��(�9�?u��LT�?.�S�̮�?l�l��?�I��I��?/�袋.�?F]t�E�?�q�q�?�q�q�?�?�?      �?                      �?              �?      �?      �?              �?      �?        ZZZZZZ�?iiiiii�?              �?�Q����?)\���(�?333333�?ffffff�?      �?      �?      �?                      �?              �?wwwwww�?�?      �?        ]t�E]�?F]t�E�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?Ց&��?����g?�?�|����?�S�n�?��8��8�?�q�q�?_�_��?�A�A�?      �?              �?      �?      �?                      �?              �?��k(��?�k(���?      �?        {�G�z�?��(\���?Y�B��?zӛ����?�$I�$I�?n۶m۶�?              �?      �?        r�q��?�q�q�?              �?      �?              �?        j�;v5,�?��"NT��?�c�1��?�s�9��?�������?�������?]t�E�?t�E]t�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?r�q��?�$I�$I�?۶m۶m�?      �?                      �?              �?n۶m۶�?�$I�$I�?      �?              �?      �?GX�i���?�{a���?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ��rD���?�и[�?e�kBP��?�	A����?�Z��D�?��4��g�?�������?������y?      �?        :�&oe�?�x+�R�?      �?      �?              �?      �?              �?        �������?�������?      �?        �������?333333�?              �?      �?        �������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?�x���!�?�C��o�?J��yJ�?�־a��?���L�?�u�)�Y�?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?�������?333333�?      �?                      �?      �?                      �?;�;��?;�;��?���Q��?)\���(�?      �?      �?UUUUUU�?�������?      �?                      �?      �?                      �?      �?        XG��).�?��:��?�rS�<��?���e�+�?      �?      �?              �?�������?�?�������?�������?      �?                      �?      �?        �?�?      �?      �?�?<<<<<<�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        ���̞?��g	�?�$I�$I�?۶m۶m�?      �?                      �?�5�5�?�Qv�Qv�?              �?W�+�ɥ?��F}g��?              �?      �?              �?        �����?��	��	�?|�W|�W�?�A�A�?      �?        �z�G��?{�G�z�?UUUUUU�?UUUUUU�?      �?                      �?�k(���?(�����?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?        �������?333333�?�rO#,��?|a���?z��y���?�a�a�?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�q�q�?              �?�?�?      �?        �������?�������?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�����?������?�������?�������?              �?      �?        r�q��?�8��8��?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?]t�E�?t�E]t�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��wrhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�=         �       
             �?�lb���?<           ��@              S                   �a@@�4���?J           P�@                                  �?l��\��?�            `w@                                   �?և���X�?             E@              
                    �?
j*D>�?             :@                                  �?      �?             (@        ������������������������       �                     @               	                   �`@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @                                   @؇���X�?             ,@                                 �Z@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                  �u@     ��?             0@                                 p`@�r����?
             .@                      	             �?����X�?             @                                   �I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?               $                   i@�5��^�?�            �t@               !                    �Q@ g�yB�?W             `@                      
             �? >��@�?U            @_@                      	          033�?      �?             0@                                   @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �        I            @[@        "       #                   @]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        %       &                   �Q@�s��=��?y            `i@        ������������������������       �                     �?        '       N                   �c@(a��䛼?x            @i@       (       ?       	          ����?H�_�r�?i            `f@        )       2                   �_@�����H�?              K@        *       1                    �?h�����?             <@       +       ,                   �]@      �?             0@        ������������������������       �                     @        -       .       	             �?ףp=
�?             $@       ������������������������       �                     @        /       0                   `Y@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        3       >                   a@���B���?             :@       4       5                    `@�J�4�?             9@        ������������������������       �                     �?        6       =                   0a@      �?             8@       7       8                   �j@z�G�z�?	             .@        ������������������������       �                      @        9       :                    �?$�q-�?             *@       ������������������������       �                     $@        ;       <                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        @       E                    \@��v��?I            @_@        A       D                    �?�<ݚ�?             "@       B       C                   Pk@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        F       G                   8p@@m���?D             ]@       ������������������������       �        '            �N@        H       M                    �? �Jj�G�?            �K@       I       L                    �J@�(\����?             D@        J       K                    �?�C��2(�?	             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �                     .@        O       P                     Q@�LQ�1	�?             7@       ������������������������       �                     2@        Q       R                   �[@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        T       �                   �f@b��H���?b            �b@       U       �                   pb@:�.���?^            �a@       V       W                    @D@�o�Nm��?O            @]@        ������������������������       �        	             *@        X       a                    �?l���B��?F             Z@        Y       \                    �K@     ��?             @@       Z       [                    �?P���Q�?             4@       ������������������������       �        
             3@        ������������������������       �                     �?        ]       ^       	          033�?r�q��?             (@       ������������������������       �                     "@        _       `                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        b                           �?*O���?4             R@       c       v                   0o@�`���?#            �H@       d       e                   �Z@���Q��?            �A@        ������������������������       �                     @        f       m                    �K@��S���?             >@       g       h                    �?����X�?             ,@        ������������������������       �                     @        i       l                    �F@�C��2(�?	             &@        j       k       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        n       s                    �M@      �?             0@       o       r                    �L@r�q��?             (@       p       q                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        t       u                   �^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        w       ~                   @f@d}h���?             ,@       x       y                   �b@8�Z$���?             *@       ������������������������       �                     @        z       {       
             �?�q�q�?             @        ������������������������       �                     �?        |       }                     K@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?���}<S�?             7@       ������������������������       �        
             .@        �       �                     N@      �?              @       ������������������������       �                     @        �       �                   p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                      @        �       �                   @E@r�q��?�            �x@        �       �       	          �����v�2t5�?            �D@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   `@�q�q�?            �@@        �       �                   �]@      �?
             0@        �       �       	          ����?      �?              @        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	          033@j���� �?             1@       �       �                     M@�q�q�?	             .@       �       �                    �?r�q��?             @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        �       �       	          ����?ȝѡ;��?�            0v@       �       �                    �R@<�U?s�?�            �r@       �       �                   h@8d[��?�            �r@       �       �                    �L@h�Y���?�            Pr@       �       �                   `\@pNho&,�?�            �n@        �       �                   �Z@���H��?             E@        ������������������������       �        
             ,@        �       �                    �?�>4և��?             <@        ������������������������       �                     @        �       �                    �?��<b���?             7@       �       �                    �?      �?             4@        �       �                   pn@      �?             @       �       �                    @I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   0n@      �?
             0@       ������������������������       �                     "@        �       �                   �n@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �o@`��7�ѝ?v            `i@       ������������������������       �        Q            �b@        �       �                    �?�1�`jg�?%            �K@        �       �                    �?z�G�z�?             $@        �       �                   �c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����?�?            �F@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                    �?     ��?              H@        �       �                    @N@���!pc�?             6@        �       �                   �]@�8��8��?             (@        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   ps@      �?             $@       �       �                   a@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �b@ȵHPS!�?             :@       �       �                   `_@�}�+r��?             3@        �       �                    @      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                    �?����X�?             @        ������������������������       �                     �?        �       �                     O@r�q��?             @        ������������������������       �                     @        �       �                    s@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?X�Cc�?$             L@        ������������������������       �                     2@        �       �                   �\@�\��N��?             C@        ������������������������       �                     @        �       �                   `c@��.k���?             A@       �       �                    �L@�g�y��?             ?@       �       �                    �?���|���?             6@        �       �                   0m@�z�G��?             $@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�8��8��?             (@       �       �                    �I@      �?              @        �       �                     G@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          033�?�����H�?             "@        �       �       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �y�@$�?�4æ�m�?��v��?=ZT"���?�������?------�?۶m۶m�?�$I�$I�?b'vb'v�?;�;��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?              �?      �?�?�������?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        o4u~�!�?��(��?����?�����?����Mb�?X9��v��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?      �?                      �?�)���d�?�Z(�c��?      �?        �F�tj�?��~�X�?���X6��?Fu�d�?�q�q�?�q�q�?�$I�$I�?�m۶m��?      �?      �?              �?�������?�������?              �?      �?      �?              �?      �?                      �?ى�؉��?��؉���?{�G�z�?�z�G��?      �?              �?      �?�������?�������?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �~j�t��?�Zd;�?�q�q�?9��8���?�$I�$I�?�m۶m��?      �?                      �?              �?�{a���?�{a��?              �?��)A��?k߰�k�?�������?333333�?F]t�E�?]t�E�?              �?      �?                      �?              �?Y�B��?��Moz��?              �?333333�?�������?              �?      �?        �|����?�����?�W|�W|�?�A�A�?Z��Y���?S2%S2%�?              �?�N��N��?�؉�؉�?      �?      �?ffffff�?�������?      �?                      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?�q�q�?և���X�?����S�?333333�?�������?      �?        �?�������?�$I�$I�?�m۶m��?      �?        F]t�E�?]t�E�?      �?      �?      �?                      �?              �?      �?      �?�������?UUUUUU�?333333�?�������?              �?      �?              �?              �?      �?      �?                      �?۶m۶m�?I�$I�$�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?        d!Y�B�?ӛ���7�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?UUUUUU�?�ڕ�]��?��+Q��?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?      �?      �?                      �?              �?              �?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�S>�6�?�b��I�?��m�>��?�C��ֲ?#�u�)��?�S�n�?�)=�$�?d�n-ܴ�?$�=����?ȝ%�淠?�0�0�?��y��y�?      �?        �$I�$I�?�m۶m��?      �?        ��,d!�?��Moz��?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?        �m۶m��?�$I�$I�?              �?      �?              �?        C���?J��8D�?      �?        A��)A�?�־a�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ��I��I�?l�l��?�������?UUUUUU�?      �?                      �?      �?              �?      �?F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?�m۶m��?�$I�$I�?      �?                      �?              �?��N��N�?�؉�؉�?�5��P�?(�����?      �?      �?      �?                      �?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?%I�$I��?�m۶m��?      �?        �5��P�?y�5���?              �?�������?�?��{���?�B!��?]t�E]�?F]t�E�?333333�?ffffff�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?      �?              �?        �q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���"hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK�h��B�<         �       
             �?�s����?F           ��@              M                    �?Ƃ<����?V           Ѐ@                                   �?��Eac��?�             k@               	       	          ����?� �	��?             I@                                    G@"pc�
�?             &@                                  @c@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        
                           �?�q�q�?            �C@                                  �K@��R[s�?            �A@                                 �g@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �                     1@                                  Pm@     ��?
             0@                                  �`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?���Q��?             $@                                  b@      �?             @        ������������������������       �                     @        ������������������������       �                     @                                  `X@      �?             @        ������������������������       �                      @                                   @L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               L                   0f@��y�+�?i            �d@              +                    �?��ۭ���?d            �c@                       
             �?d��0u��?             >@        ������������������������       �                     @        !       *                   xr@�+e�X�?             9@       "       '                   �c@�q�q�?             8@       #       &                   �N@�X�<ݺ?             2@        $       %                    `Q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        (       )       	          ���@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ,       7                    �K@��7PB��?O            �_@       -       .                   ``@p�|�i�?-             S@        ������������������������       �                    �@@        /       6       	          ����?Du9iH��?            �E@       0       5       	          ����?     ��?             @@       1       2                   �`@`Jj��?             ?@       ������������������������       �                     9@        3       4                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        8       E                   0b@t�F�}�?"            �I@       9       D                   @x@(N:!���?            �A@       :       C                    `@l��\��?             A@       ;       B                   �`@H%u��?             9@        <       A                    �?���!pc�?
             &@       =       @                   �_@z�G�z�?	             $@       >       ?       
             �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �                     "@        ������������������������       �                     �?        F       G       	          833�?      �?             0@        ������������������������       �                     @        H       K                    �?�θ�?             *@       I       J                   �b@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        N                           �?Ї	{�k�?�             t@       O       P                   �U@|)����?�            q@        ������������������������       �                      @        Q       x       	          `ff @�3ظ\�?�            �p@       R       m                   �b@P�19A'�?�             j@       S       T                   �e@`ۘV�?j            @e@        ������������������������       �        $            �K@        U       V                   �f@d����?F            �\@        ������������������������       �                      @        W       X                    �F@h��)�~�?E            @\@        ������������������������       �        
             1@        Y       `                    @G@��8����?;             X@        Z       [                   �`@���Q��?             $@        ������������������������       �                     @        \       ]                    �?z�G�z�?             @        ������������������������       �                      @        ^       _       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        a       l                   (q@����"$�?5            �U@       b       c                    @L@�^����?"            �M@        ������������������������       �                     8@        d       e                   �Z@z�G�z�?            �A@        ������������������������       �                     @        f       k                    �M@��a�n`�?             ?@        g       j                    q@�z�G��?             $@       h       i                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             5@        ������������������������       �                     ;@        n       w                    �Q@:�&���?            �C@       o       r                    �?�#-���?            �A@        p       q                    �H@      �?              @        ������������������������       �                      @        ������������������������       �                     @        s       v                   �b@ 7���B�?             ;@        t       u                    @H@�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     0@        ������������������������       �                     @        y       ~                    j@�g�y��?&             O@        z       {                   @b@���}<S�?             7@       ������������������������       �                     3@        |       }       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �C@        �       �                   �`@ \� ���?"            �H@       �       �                   �Y@�X�<ݺ?             B@        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?XB���?             =@       �       �                     N@P���Q�?             4@        �       �                   @^@�����H�?             "@        �       �                    `@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     "@        �       �       	          @33�?�θ�?	             *@        ������������������������       �                     �?        �       �       	          `ff�?r�q��?             (@       �       �                   �l@�C��2(�?             &@       ������������������������       �                     @        �       �       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?Xf�?s��?�            �w@       �       �       	          `ff @�É`��?�            �t@       �       �                    �?$΅9>��?�            `t@        �       �                   �_@������?;             \@        �       �                    �I@� �	��?             I@       �       �                   i@П[;U��?             =@        �       �                    �?d}h���?             ,@        ������������������������       �                     �?        �       �                    �?8�Z$���?             *@       ������������������������       �                     @        �       �                    @D@      �?              @        ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?�r����?	             .@       �       �       	          ����?�C��2(�?             &@       �       �                    @F@ףp=
�?             $@        �       �                   �q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �o@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@����X�?             5@       �       �                   `a@և���X�?             @       �       �                    \@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   Pj@؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        �       �                   �b@�חF�P�?             O@       �       �       	          ����?4և����?             L@       �       �                    @N@�X�<ݺ?             K@       ������������������������       �                    �I@        ������������������������       �                     @        ������������������������       �                      @        �       �                    �J@r�q��?             @       �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?Xφ���?�            �j@        �       �                    c@6YE�t�?            �@@       �       �                    �G@ 	��p�?             =@        ������������������������       �                     $@        �       �                   �f@�KM�]�?             3@        ������������������������       �                     �?        �       �                   0s@�X�<ݺ?             2@       ������������������������       �                     .@        �       �                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �O@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �S@0m��5!�?z            �f@        �       �                    @�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                   @n@��f�{��?t            �e@       ������������������������       �        ?             X@        �       �                   @[@P�Lt�<�?5             S@        �       �                   @q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    _@`׀�:M�?3            �R@        �       �       	          @33�?�nkK�?             7@       ������������������������       �                     3@        �       �                   �^@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �I@        ������������������������       �                      @        �       �                    �G@      �?             G@        �       �                    �?�θ�?             *@        �       �                    �F@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �J@����e��?            �@@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�q�����?             9@       �       �                   Pd@@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �                     &@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ��mQ��?-I׺��?�e���?��U���?&���^B�?�%���^�?�Q����?)\���(�?F]t�E�?/�袋.�?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?X|�W|��?PuPu�?�k(���?(�����?              �?      �?              �?      �?�������?UUUUUU�?      �?                      �?�������?333333�?      �?      �?      �?                      �?      �?      �?              �?      �?      �?              �?      �?                      �?�������?�ˊ���?�Kz���?�?m�K�?wwwwww�?DDDDDD�?      �?        ���Q��?R���Q�?�������?UUUUUU�?�q�q�?��8��8�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        I$�D"�?�v��n��?^Cy�5�?�k(����?              �?w�qGܱ?qG�w��?      �?      �?�B!��?���{��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?777777�?�A�A�?|�W|�W�?�������?------�?���Q��?)\���(�?t�E]t�?F]t�E�?�������?�������?�q�q�?�q�q�?      �?                      �?      �?              �?                      �?              �?      �?              �?      �?              �?ى�؉��?�؉�؉�?      �?      �?      �?                      �?      �?              �?        �O���?6�l�?h�h��?��/��/�?      �?        /R�Dȴ?���f�?<�7c�?,���?�������?�������?              �?�(�j�?�����a�?      �?        Ź�Q��?�(�u���?              �?UUUUUU�?UUUUUU�?�������?333333�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        6eMYSִ?YS֔5e�?W'u_�?u_[4�?              �?�������?�������?      �?        �c�1Ƹ?�s�9��?333333�?ffffff�?      �?      �?      �?                      �?      �?                      �?              �?�o��o��?�A�A�?_�_�?�A�A�?      �?      �?      �?                      �?h/�����?	�%����?F]t�E�?]t�E�?      �?                      �?              �?      �?        �B!��?��{���?d!Y�B�?ӛ���7�?              �?      �?      �?              �?      �?                      �?և���X�?
^N��)�?�q�q�?��8��8�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        �{a���?GX�i���?�������?ffffff�?�q�q�?�q�q�?      �?      �?              �?      �?                      �?              �?              �?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?]t�E�?F]t�E�?      �?              �?      �?      �?                      �?              �?�8�{n�?a�+F�? K���?�Ӛ��?{�r��b�?f5�8t�?I�$I�$�?n۶m۶�?)\���(�?�Q����?�{a���?��=���?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?              �?      �?      �?              �?      �?        �������?�?]t�E�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?              �?      �?        �$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?�������?333333�?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?�Zk����?��RJ)��?I�$I�$�?�m۶m۶?��8��8�?�q�q�?      �?                      �?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?���z��?�rp�_��?'�l��&�?e�M6�d�?������?�{a���?      �?        �k(���?(�����?              �?��8��8�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        kdu�J�?�rS�<��?9��8���?�q�q�?      �?                      �?������?�}A_Ї?      �?        ���k(�?(�����?      �?      �?              �?      �?        ��L��?к����?�Mozӛ�?d!Y�B�?      �?              �?      �?      �?                      �?      �?                      �?      �?      �?ى�؉��?�؉�؉�?      �?      �?              �?      �?              �?        6�d�M6�?e�M6�d�?      �?      �?      �?                      �?���Q��?�p=
ף�?�$I�$I�?n۶m۶�?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�|�PhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK�h��B�<         �       
             �?�$�����?9           ��@                                 �a@�A����?K           ��@                      	          033�?�&/�E�?S             _@                                 `X@�D�e���?;            @U@               
                   `Q@      �?
             0@                                  �?�r����?	             .@       ������������������������       �                      @               	                    V@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        1            @Q@                                  �U@�ݜ�?            �C@        ������������������������       �                      @                                  �c@�L���?            �B@       ������������������������       �                     >@                                   @M@և���X�?             @        ������������������������       �                     @                                  �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?               Q                    �?�����?�            `y@               L                    �?(Q��h�?h            @d@              %                    �?      �?T             `@               "                   �b@r�q��?             B@                     	          ����?`Jj��?             ?@        ������������������������       �                     ,@               !       	             �?�t����?             1@                                  �o@���Q��?             @        ������������������������       �                      @                                    @�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        #       $                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        &       A                   �`@nM`����?;             W@       '       :                   0p@�������?%             N@       (       )       
             �?*O���?             B@        ������������������������       �                     @        *       9                    �N@     ��?             @@       +       ,                   �\@|��?���?             ;@        ������������������������       �                     �?        -       2                    �?��
ц��?             :@        .       1                   �c@"pc�
�?             &@        /       0                    _@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        3       4                   �a@�q�q�?	             .@       ������������������������       �                      @        5       6                    @G@����X�?             @        ������������������������       �                     @        7       8       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ;       @                   �e@      �?             8@       <       =                   `r@"pc�
�?             6@       ������������������������       �                     ,@        >       ?                   `s@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        B       C       
             �?     ��?             @@        ������������������������       �                     �?        D       E                   pb@��� ��?             ?@       ������������������������       �                     1@        F       G                   �b@����X�?	             ,@        ������������������������       �                     �?        H       I                    d@�θ�?             *@       ������������������������       �                     "@        J       K                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        M       N                   �S@@�0�!��?             A@        ������������������������       �                     @        O       P                   f@��a�n`�?             ?@       ������������������������       �                     <@        ������������������������       �                     @        R       U                   �Z@�&�4rd�?�            �n@        S       T                   `n@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        V       �                   �b@� g\z�?�            �m@       W       X                   `[@py�����?�             l@        ������������������������       �                     C@        Y       d                    \@0�#�.^�?i            `g@        Z       c                    �?      �?
             0@       [       ^                     L@����X�?	             ,@        \       ]       	             �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        _       `                   Pr@�����H�?             "@       ������������������������       �                     @        a       b       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        e       l                   �[@�����?_            `e@        f       g                   `_@����X�?             ,@        ������������������������       �                     @        h       k                   �n@      �?              @       i       j                    b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        m       |                    �?�������?X            �c@        n       {                   hu@������?             >@       o       z                   `c@d}h���?             <@       p       w                    �?�����?
             3@       q       r                    �H@z�G�z�?             .@        ������������������������       �                     �?        s       t                    �?؇���X�?             ,@       ������������������������       �                     $@        u       v                    �I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        x       y       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        }       �                    �?����}��?I            �_@       ~       �                    `@ �ׁsF�?:             Y@               �       	          `ff�?@��8��?             H@        ������������������������       �                     4@        �       �                   �_@h�����?             <@       ������������������������       �                     8@        �       �                    �?      �?             @       �       �                   pk@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     J@        ������������������������       �                     ;@        �       �                    �?X�Cc�?
             ,@       �       �                   p@ףp=
�?             $@       ������������������������       �                     @        �       �       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�v�����?�            @x@        �       �                   @E@�.̦˝�?V             a@        �       �                    @M@      �?             @@       �       �                   `\@�X�<ݺ?             2@        �       �                   `^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                   �^@      �?	             ,@        ������������������������       �                     @        �       �                    �?���|���?             &@        �       �                     P@z�G�z�?             @        ������������������������       �                     @        �       �                    �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          033�?      �?             @       �       �                    [@���Q��?             @        ������������������������       �                      @        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?$+ޠ�5�?A            @Z@       �       �                   `\@:���u��?/            @S@        �       �                    �?�LQ�1	�?             7@        ������������������������       �                     @        �       �       	          tff�?      �?             4@       �       �                    �?�q�q�?	             .@       �       �                   �l@r�q��?             (@        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �       	          ����?      �?             @        ������������������������       �                     �?        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   (t@�>����?!             K@       �       �                   �j@�IєX�?            �I@        �       �                   �h@�LQ�1	�?             7@       ������������������������       �        
             3@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @J@X�Cc�?             <@        ������������������������       �                     @        �       �                   �h@�eP*L��?             6@        ������������������������       �                     @        �       �                    �L@j���� �?
             1@        �       �                    a@      �?              @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	             �?�q�q�?             "@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    @Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �g@��H�$�?�            `o@       �       �                    @h�U���?�             o@       �       �                    �?0x�!���?�            �m@        ������������������������       �        +            @R@        �       �                   �a@�6,r➷?e            �d@        �       �       	          `ff�?�8��8��?             H@       ������������������������       �                     F@        ������������������������       �                     @        �       �       	             @ȑ����?F            @]@       �       �                    c@�]���?D            �\@       �       �                    �?����r�??            �[@       ������������������������       �        "             M@        �       �                   @[@ pƵHP�?             J@        �       �                    �?      �?             @       �       �       	          ����      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     H@        �       �                    �K@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���!pc�?             &@       ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                     I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�B0  3O��k�?g���-J�?үz�@�?T�ѯz�?�s�9�?2�c�1�?�???????�?      �?      �?�?�������?              �?�$I�$I�?�m۶m��?              �?      �?                      �?              �?�i�i�?\��[���?      �?        L�Ϻ��?}���g�?              �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?�U�3���?���
�?������?x�5?,�?      �?      �?�������?UUUUUU�?���{��?�B!��?      �?        <<<<<<�?�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �������?�������?              �?      �?        zӛ����?C���,�?�������?�������?�q�q�?�q�q�?      �?              �?      �?{	�%���?	�%����?              �?�;�;�?�؉�؉�?/�袋.�?F]t�E�?333333�?�������?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?F]t�E�?/�袋.�?              �?      �?      �?      �?                      �?      �?              �?      �?      �?        �B!��?�{����?              �?�$I�$I�?�m۶m��?      �?        �؉�؉�?ى�؉��?              �?      �?      �?      �?                      �?�������?ZZZZZZ�?      �?        �c�1Ƹ?�s�9��?              �?      �?        i�>�%C�?&C��6��?333333�?�������?      �?                      �?Z����?u�c�D@�?I�7�&��?�*;L�?              �?w��?��b���?      �?      �?�$I�$I�?�m۶m��?333333�?�������?      �?                      �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        d7��Dv�?�Md7��?�$I�$I�?�m۶m��?              �?      �?      �?�������?�������?      �?                      �?              �?b��x�Y�?�fue*�?�?wwwwww�?۶m۶m�?I�$I�$�?^Cy�5�?Q^Cy��?�������?�������?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?      �?      �?                      �?              �?      �?        �@ �?����~��?{�G�z�?�G�z��?UUUUUU�?UUUUUU�?              �?�$I�$I�?�m۶m��?              �?      �?      �?      �?      �?      �?                      �?              �?              �?              �?%I�$I��?�m۶m��?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?Jd����?�n�'�i�?�[�w��?<�H��?      �?      �?�q�q�?��8��8�?      �?      �?              �?      �?                      �?      �?      �?      �?        F]t�E�?]t�E]�?�������?�������?              �?      �?      �?      �?                      �?      �?      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �K��K��?�h��h��?dj`��?qV~B���?d!Y�B�?Nozӛ��?      �?              �?      �?UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?�������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�Kh/��?h/�����?�?�?��Moz��?Y�B��?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?%I�$I��?              �?]t�E�?t�E]t�?              �?�������?ZZZZZZ�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�$Ԑ�W�?���򖄪?�����?��"NT��?��~���?�5�5�?      �?        s�,��r�?�0�Ө?UUUUUU�?UUUUUU�?      �?                      �?��~���?���?��ʇq�?���ϑ?�oX����?��)A��?      �?        'vb'vb�?;�;��?      �?      �?      �?      �?      �?                      �?      �?              �?        �������?�������?      �?                      �?              �?F]t�E�?t�E]t�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ6pWAhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM)hzh)h,K ��h.��R�(KM)��h��B@J         �                    �?��t�?:           ��@              =       	          ����?l�:���?0           @               *                    �?�0u��A�?m            �f@                                 ``@0˚p&��?A            @[@                                   �?��|�5��?            �G@                                  @[@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        	              
             �?�����H�?             B@       
              	             �? 7���B�?             ;@       ������������������������       �                     :@        ������������������������       �                     �?                                   X@�q�q�?             "@        ������������������������       �                     @                                  @`@      �?             @                                 �X@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                  @E@Z��Yo��?$             O@        ������������������������       �                     $@                                  �b@      �?             J@                                  �x@`2U0*��?             9@       ������������������������       �        
             8@        ������������������������       �                     �?               !                    n@X�<ݚ�?             ;@                                   �\@d}h���?             ,@                                   �?      �?             @        ������������������������       �                      @                                  �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        "       '                   �r@�	j*D�?
             *@       #       $                   p`@�����H�?             "@       ������������������������       �                     @        %       &                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        (       )                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        +       6                   �b@���BK�?,            �Q@       ,       -                   �j@Ԫ2��?$            �L@       ������������������������       �                     @@        .       3       
             �?`�Q��?             9@       /       2                    \@�����H�?             2@        0       1       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             .@        4       5                    �H@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        7       8                    h@d}h���?             ,@        ������������������������       �                     �?        9       <                   Pd@8�Z$���?             *@       :       ;                   �c@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        >       ?                   �U@��10��?�            �s@        ������������������������       �                      @        @       {       
             �?��K]�?�            �s@       A       R                    �?�E�J��?�            �p@        B       Q                    �?����X�?            �A@       C       P                    �?J�8���?             =@       D       K                   �`@l��
I��?             ;@        E       F                    �G@      �?             (@        ������������������������       �                     @        G       J                     L@؇���X�?             @        H       I       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        L       M                   �u@�r����?
             .@       ������������������������       �                     &@        N       O                   pc@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        S       l                   �`@@\�*��?�            @m@        T       Y                    @J@b �57�?@            �Y@        U       V                    a@@��8��?             H@       ������������������������       �                    �D@        W       X                   �a@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        Z       [                   @R@lGts��?'            �K@        ������������������������       �                     �?        \       e                    \@h�WH��?&             K@        ]       b       	             @������?             1@       ^       _                    @L@؇���X�?	             ,@        ������������������������       �                     @        `       a                    �L@      �?              @        ������������������������       �                      @        ������������������������       �                     @        c       d                   �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        f       k                    �L@�?�|�?            �B@        g       j                   �\@@4և���?             ,@        h       i       	             @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             (@        ������������������������       �                     7@        m       t                   q@�z�N��?O            ``@       n       o                   �_@�K}��?:            �Y@       ������������������������       �        &            �P@        p       s                   `@������?             B@        q       r                    �F@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ?@        u       x                    c@ 	��p�?             =@       v       w                    �Q@ 7���B�?             ;@       ������������������������       �                     :@        ������������������������       �                     �?        y       z                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        |       �       	          033�?��+7��?             G@        }       ~                    @D@      �?
             0@        ������������������������       �                      @               �                    �?և���X�?	             ,@       �       �                     J@�eP*L��?             &@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@�r����?             >@       �       �       	          `ff @ܷ��?��?             =@       �       �                    @N@؇���X�?             5@       �       �                   @`@      �?             (@        ������������������������       �                     @        �       �                   �^@և���X�?             @        ������������������������       �                      @        �       �                    �?z�G�z�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?���w~��?
           Pz@       �       �                   �`@��ED���?�             p@        �       �       	          �����{ /h��?3            �S@        ������������������������       �                     @        �       �                   `T@�E����?1             R@        �       �       
             �?     ��?             0@       �       �                    @K@@4և���?
             ,@        ������������������������       �                     @        �       �                   �X@      �?              @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   Pt@�>4և��?%             L@       �       �                    �L@���c���?"             J@        �       �                    �?h�����?             <@       ������������������������       �                     ;@        ������������������������       �                     �?        �       �                    @M@      �?             8@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��s����?             5@        ������������������������       �                     &@        �       �       
             �?���Q��?             $@        �       �                    �?      �?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?r�q��?             @        �       �                    \@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �O@�IQu`�?r            �f@        �       �                   @_@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �q@XpBt,��?o            �e@       �       �       	          pff�?�?�|�?\            �b@       �       �                    �?`Ql�R�?W            �a@       �       �                   �[@`o��b�?L             _@        �       �                   �o@��S�ۿ?	             .@       ������������������������       �                     (@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        C            @[@        �       �                   �m@�t����?             1@       ������������������������       �                     &@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   l@؇���X�?             @        ������������������������       �                     @        �       �                   Pn@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@�+$�jP�?             ;@        �       �                   �b@      �?             $@        ������������������������       �                     @        �       �                    �?����X�?             @        �       �                   �s@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@        �                          �?B\Q���?e            `d@       �       �                    �?&RN���?A            @Z@        �       �                   `X@     ��?             @@        ������������������������       �                      @        �       �       	          ����?(;L]n�?             >@        �       �                    �?�C��2(�?             &@       �       �                    q@؇���X�?             @       ������������������������       �                     @        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             3@        �                          �?P�t��?.            @R@       �       �                    �F@x�K��?             �I@        �       �                    �?؇���X�?             @        �       �                     D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �             	          `ff�?�X����?             F@       �                          �P@      �?             :@       �       �                    �?\X��t�?             7@        �       �       	          pff�?r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �                    N@���!pc�?
             &@        ������������������������       �                     �?        �       �       	          ����?z�G�z�?	             $@        ������������������������       �                     �?        �             	          ����?�����H�?             "@                                  d@      �?             @        ������������������������       �                      @                                �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              
                  @a@�X�<ݺ?	             2@              	                  �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     0@                    
             �?8�A�0��?             6@                                 O@��.k���?
             1@                   	          ����?���|���?             &@        ������������������������       �                     @                                 _@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                 @r�q��?             @        ������������������������       �                     @                    
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 _@J�8���?$             M@        ������������������������       �                     4@              "                  �l@�\��N��?             C@                               �`@�GN�z�?             6@                                �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @               !                   �?      �?	             0@       ������������������������       �                     .@        ������������������������       �                     �?        #      $                  �m@     ��?             0@        ������������������������       �                     @        %      &                   o@�z�G��?             $@        ������������������������       �                      @        '      (                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM)KK��hb�B�  |&�{&��?�l�l�?�%'��?�6�B^�?�������?�������?����[�?#s�3R�?x6�;��?br1���?]t�E]�?F]t�E�?              �?      �?        �q�q�?�q�q�?h/�����?	�%����?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?      �?              �?      �?              �?        !�B!�?���{��?              �?      �?      �?���Q��?{�G�z�?      �?                      �?r�q��?�q�q�?I�$I�$�?۶m۶m�?      �?      �?              �?      �?      �?              �?      �?              �?        ;�;��?vb'vb'�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?      �?              �?      �?        $Zas �?��RO�o�?p�}��?$���>��?              �?{�G�z�?��(\���?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?        I�$I�$�?۶m۶m�?              �?;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��u�?*���\��?      �?        ���?�˿�˿�?��~���?�-���?�$I�$I�?�m۶m��?|a���?�rO#,��?h/�����?Lh/����?      �?      �?              �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?        �?�������?              �?      �?      �?              �?      �?              �?                      �?^�^�?���?�H%�e�?��VC��?UUUUUU�?UUUUUU�?              �?�$I�$I�?۶m۶m�?      �?                      �?�־a�?�<%�S��?      �?        B{	�%��?��^B{	�?�?xxxxxx�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?к����?*�Y7�"�?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?              �?ձ�6Ls�?qBJ�eD�?�?�������?              �?�q�q�?�q�q�?�������?�������?      �?                      �?              �?�{a���?������?h/�����?	�%����?              �?      �?              �?      �?      �?                      �?Y�B��?zӛ����?      �?      �?      �?        ۶m۶m�?�$I�$I�?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�?�������?a���{�?��=���?�$I�$I�?۶m۶m�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?              �?      �?        ۸�*��?J�ު� �?�'�	�?��=aO��?�A�A�?�|˷|��?              �?r�q��?�q�q�?      �?      �?�$I�$I�?n۶m۶�?              �?      �?      �?      �?      �?      �?                      �?              �?      �?        �$I�$I�?�m۶m��?;�;��?�;�;�?�m۶m��?�$I�$I�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?z��y���?�a�a�?      �?        333333�?�������?      �?      �?      �?      �?              �?      �?                      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?              �?�`�`�?��I��I�?333333�?�������?      �?                      �?L�w�Z�?�>���T�?*�Y7�"�?к����?}g���Q�?W�+�ɕ?���{��?�B!��?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        <<<<<<�?�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        /�����?B{	�%��?      �?      �?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ���A2��?/����?�����?]ʥ\ʥ�?      �?      �?              �?�������?�?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?              �?        ˖-[�l�?�4iҤI�?�?ssssss�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        ]t�E]�?�E]t��?      �?      �?��Moz��?!Y�B�?UUUUUU�?�������?      �?                      �?F]t�E�?t�E]t�?              �?�������?�������?              �?�q�q�?�q�q�?      �?      �?      �?              �?      �?              �?      �?              �?              �?        �q�q�?��8��8�?      �?      �?              �?      �?                      �?/�袋.�?颋.���?�������?�?F]t�E�?]t�E]�?      �?              �?      �?      �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?|a���?�rO#,��?              �?y�5���?�5��P�?�袋.��?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?      �?              �?333333�?ffffff�?      �?              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ2��JhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@A         �                    �?��/.��?N           ��@              ;       	          ����?4`�/Z�?=           P@                      
             �?���r
��?y            @h@                                 �_@�(�,�J�?C            �]@                     	          ����?�.ߴ#�?"            �N@       ������������������������       �        !             M@        ������������������������       �                     @                      	          833�?��h!��?!            �L@       	       
                   �b@ >�֕�?            �A@       ������������������������       �                     ?@                                   �G@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   b@���|���?
             6@                                 �g@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     @                                  `X@      �?6             S@        ������������������������       �                     @               ,                    �?��oh���?5            @R@                                  �E@X�;�^o�?(            �K@                                   @C@����X�?	             ,@        ������������������������       �                     @                                   @D@X�<ݚ�?             "@        ������������������������       �                      @                                  �c@����X�?             @                                 �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                %                    �?��p\�?            �D@        !       $       	          @33�?�����H�?             "@       "       #                   �d@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        &       '                   �^@      �?             @@        ������������������������       �        	             .@        (       +                   `d@�t����?             1@       )       *                    �M@      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �                     �?        -       8                    �?      �?             2@       .       3                    b@և���X�?
             ,@        /       0                    �?r�q��?             @        ������������������������       �                     @        1       2                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        4       7                   �d@      �?              @       5       6                    �N@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        9       :                   @b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        <       �                   �u@0-�Z��?�            0s@       =       >                   �U@��5�l@�?�            Pr@        ������������������������       �                      @        ?       z       
             �?��_F	��?�            0r@       @       w                    `R@���N8�?�            �o@       A       b                   P`@���i��?�            @o@        B       Q                    �?0{�v��?K            @_@       C       J                   �r@@9G��?9            �X@       D       I                   @Z@�|���?4             V@        E       F                    �L@$�q-�?             *@       ������������������������       �                     "@        G       H                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        ,            �R@        K       L                    s@�z�G��?             $@        ������������������������       �                      @        M       P                    @I@      �?              @        N       O                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        R       a       	          ����?�+$�jP�?             ;@       S       ^                   �q@�t����?             1@       T       ]       	          ����?d}h���?	             ,@       U       V                   �]@8�Z$���?             *@        ������������������������       �                     �?        W       X                    `@�8��8��?             (@        ������������������������       �                     @        Y       \                    @M@      �?              @        Z       [                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        _       `                    @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        c       d                    �?@�n�1�?R            @_@        ������������������������       �                     =@        e       v                   �b@@��8��??             X@       f       i                    �D@���#�İ?+            �M@        g       h                    �C@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        j       k                    �?�h����?(             L@        ������������������������       �                     @        l       u                    �?p���?#             I@       m       t                   �a@г�wY;�?             A@       n       o                     M@P���Q�?             4@       ������������������������       �        
             $@        p       s                    @N@ףp=
�?             $@        q       r       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             ,@        ������������������������       �        
             0@        ������������������������       �                    �B@        x       y                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        {       �       	          033@��Sݭg�?            �C@       |       }                    �?�'�`d�?            �@@        ������������������������       �                      @        ~       �                    c@�חF�P�?             ?@              �                    @N@$�q-�?             :@       �       �                    @J@؇���X�?             ,@        ������������������������       �                     @        �       �       	          `ff�?�<ݚ�?             "@       �       �                   Pm@      �?              @       ������������������������       �                     @        �       �                    c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?և���X�?             ,@        �       �                   �_@      �?              @        ������������������������       �                     �?        �       �                     L@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��91��?           z@       �       �                    �K@�n����?�            �u@       �       �       	          ����?<I����?�            �n@       �       �                   �`@���{h�?�            `l@        �       �                    @�����H�?             B@       �       �       
             �?�#-���?            �A@        �       �                   �v@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @c@�g�y��?             ?@        ������������������������       �                     �?        ������������������������       �                     >@        ������������������������       �                     �?        �       �                   �c@�X�T���?w            �g@        �       �                   �b@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �a@@i�)ԙ�?q            �f@        �       �       
             �? ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@        �       �                   @^@�(�Tw�?d            �c@        �       �                    @E@г�wY;�?+             Q@        ������������������������       �                     C@        �       �                    �H@��S�ۿ?             >@       �       �                    \@      �?             0@        ������������������������       �                     @        �       �                   �p@z�G�z�?	             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             ,@        ������������������������       �        9             V@        �       �       
             �?p�ݯ��?
             3@       �       �                    �?      �?             0@        ������������������������       �                     @        �       �                     I@$�q-�?             *@       ������������������������       �                     $@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @O@
�c�Z�?F             Y@       �       �                   �O@�q�q�?,             N@        ������������������������       �                      @        �       �                   �h@θ	j*�?&             J@        ������������������������       �                      @        �       �                   �m@�zv�X�?              F@       �       �                   `_@և���X�?             5@        ������������������������       �                     @        �       �                    �L@      �?             0@        ������������������������       �                     @        �       �                   pb@���Q��?
             $@        �       �                   @e@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���Q��?             @       �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �_@��<b���?             7@        �       �                    �?      �?             @       �       �       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @L@�KM�]�?             3@        �       �                    �?�q�q�?             @        ������������������������       �                      @        �       �       	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        �       �                    �?ףp=
�?             D@       �       �       	          ����?��S�ۿ?             >@        �       �                   (s@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     6@        �       �       	          ����?z�G�z�?             $@        ������������������������       �                     @        �       �       	          ���@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �J@^|�_��?0            �Q@        �       �                    �?¦	^_�?             ?@        ������������������������       �                      @        �       �                   �c@�û��|�?             7@        ������������������������       �                     @        �       �       	          ����?�d�����?	             3@       ������������������������       �                     (@        �       �       
             �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?�z�G��?             D@        �       �       
             �?X�<ݚ�?             2@       �       �                    @N@�q�q�?	             (@        �       �                   �`@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �                         �j@�C��2(�?             6@        �                          @�<ݚ�?	             "@       �                          �?      �?              @                                  �M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        �t�bh�h)h,K ��h.��R�(KMKK��hb�BP  �"�Zw�?6�n�R��?���9��?V��1�:�?���fy�?�<�L�v�?_[4��?h8�����?XG��).�?�K�`m�?              �?      �?        p�}��?Hp�}�?�A�A�?��+��+�?              �?      �?      �?      �?                      �?]t�E]�?F]t�E�?�������?�?              �?      �?                      �?      �?      �?              �?ȏ?~��?����?�־a��?J��yJ�?�m۶m��?�$I�$I�?      �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �]�ڕ��?��+Q��?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?      �?      �?        <<<<<<�?�?      �?      �?      �?                      �?              �?      �?      �?�$I�$I�?۶m۶m�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?�������?              �?      �?              �?              �?      �?              �?      �?        =m�\+�?Xn�z��?(���"��?�b���`�?      �?        P��Z�?>�m���?�a�a�?��y��y�?�I+��?d;�O���?;�O��n�?V-��?9/���?������?F]t�E�?��.���?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?              �?333333�?ffffff�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?B{	�%��?/�����?�������?�������?۶m۶m�?I�$I�$�?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?����Mb�?�rh��|�?              �?UUUUUU�?UUUUUU�?'u_[�?��N��?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?{�G�z�?\���(\�?�?�?�������?ffffff�?              �?�������?�������?      �?      �?              �?      �?                      �?              �?              �?              �?      �?      �?              �?      �?        �i�i�?�|˷|��?'�l��&�?6�d�M6�?      �?        ��RJ)��?�Zk����?;�;��?�؉�؉�?�$I�$I�?۶m۶m�?              �?�q�q�?9��8���?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?333333�?�������?      �?                      �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?                      �?��Յf�?����e�?��L|�w�?F5�� �?f�_��e�?�M!д?�9�K��?��gG�?�q�q�?�q�q�?�A�A�?_�_�?      �?      �?      �?                      �?��{���?�B!��?              �?      �?                      �?�|�pT�?:kP<�q�?�q�q�?�q�q�?      �?                      �?��x��x�?��?O��N���?;�;��?              �?      �?        p��o���?�A�A�?�?�?      �?        �������?�?      �?      �?      �?        �������?�������?      �?                      �?      �?              �?        Cy�5��?^Cy�5�?      �?      �?      �?        ;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        ���Q��?���(\��?�������?�������?              �?�؉�؉�?�N��N��?      �?        ��.���?�袋.��?۶m۶m�?�$I�$I�?      �?              �?      �?              �?�������?333333�?�������?�������?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ��,d!�?��Moz��?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�k(���?(�����?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        �������?�������?�������?�?      �?      �?      �?                      �?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �ԓ�ۥ�?�6��?��Zk���?�RJ)���?      �?        8��Moz�?��,d!�?              �?Cy�5��?y�5���?      �?        �$I�$I�?�m۶m��?              �?      �?        333333�?ffffff�?r�q��?�q�q�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        F]t�E�?]t�E�?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�phG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�D         �                    �?���ƒ�?C           ��@              �       	          033�?���t���?T           H�@                                 @E@�r�؜�?-           P~@               	       
             �?����?�?1            @T@                                  �?�]0��<�?"            �N@       ������������������������       �                     H@                      
             �?8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        
                           �?�G�z��?             4@                                 �a@���Q��?             $@                                 �\@�q�q�?             "@                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                      	          ����?�z�G��?             $@                                  �?      �?              @                                  `_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @               l       	             �?h#E�Y�?�            @y@              C       
             �?fP*L��?�            @s@               0                   `m@     ��?'             P@                                 �_@h+�v:�?             A@        ������������������������       �                     @                                   �?�c�Α�?             =@        ������������������������       �                     $@                )                   k@D�n�3�?             3@       !       (                   0a@�<ݚ�?             "@       "       '                    �K@�q�q�?             @       #       $                   �g@�q�q�?             @        ������������������������       �                     �?        %       &                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        *       /       	          ����?ףp=
�?             $@       +       ,                    �?�q�q�?             @        ������������������������       �                     �?        -       .                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        1       :                   �p@�������?             >@        2       3                   �_@      �?             0@        ������������������������       �                     @        4       9                   �`@"pc�
�?             &@        5       6                    �?�q�q�?             @        ������������������������       �                     @        7       8                   po@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ;       B                    �?X�Cc�?	             ,@        <       =       	          ����?����X�?             @        ������������������������       �                      @        >       ?                    �?���Q��?             @        ������������������������       �                      @        @       A                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        D       Y                    �?p��Gӹ?�            �n@        E       L                    �?:	��ʵ�?"            �F@        F       K                   @]@և���X�?             ,@        G       H                    @I@؇���X�?             @        ������������������������       �                     @        I       J                   �k@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        M       N                   �k@`Jj��?             ?@        ������������������������       �                     .@        O       X       	          ����?      �?             0@       P       Q                    �?؇���X�?             ,@        ������������������������       �                     @        R       W                   �b@"pc�
�?
             &@       S       V                    ]@ףp=
�?	             $@        T       U                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        Z       k                   0h@��}�
�?}            �h@       [       j                   �d@��F�D�?|            �h@       \       g                   pd@ ��+,��?O            @_@       ]       ^                    @L@p�,�V��?M            @^@       ������������������������       �        <            @X@        _       f                   �s@�8��8��?             8@       `       e                    �?�nkK�?             7@        a       d                    �?�����H�?             "@       b       c                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        h       i                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        -            @R@        ������������������������       �                     �?        m       x                    �?r�qG�?6             X@        n       w                   8q@l��[B��?             =@       o       v       	          ����?����X�?             5@       p       q                    �?r�q��?             2@        ������������������������       �                     �?        r       s                   �`@�t����?
             1@       ������������������������       �                     &@        t       u                    @L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        y       �                   r@� y���?&            �P@       z       �                   pq@��[�8��?            �I@       {       |                   �Z@�����H�?            �F@        ������������������������       �                      @        }       ~                   �b@Du9iH��?            �E@        ������������������������       �                     .@               �                   �\@ �Cc}�?             <@        ������������������������       �                     �?        �       �       	          033�?�>����?             ;@        �       �                    �?���Q��?             @       �       �                   @e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     @        ������������������������       �                     0@        �       �                    l@�t����?'             Q@       �       �       	          ���@r�q��?             B@       �       �       	          `ff@�θ�?             :@       �       �                   pc@"pc�
�?             6@       �       �                    @      �?
             0@       ������������������������       �        	             .@        ������������������������       �                     �?        �       �                   `T@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?     ��?             @@        �       �       	          ���@�θ�?             *@       �       �                   �]@      �?              @        ������������������������       �                     @        �       �                     J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    ]@D�n�3�?             3@        ������������������������       �                      @        �       �       	          033@ҳ�wY;�?             1@        �       �                   �d@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        �       �       	           33@�q�q�?             @       �       �                   �l@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                         �b@�I
��#�?�            �v@       �       �                    �?d#,����?�            �t@        �       �       	          033@�c�Α�?             =@       �       �                   �a@�LQ�1	�?             7@       �       �                   �j@��.k���?             1@        �       �                   �_@z�G�z�?             @        ������������������������       �                     @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?�q�q�?
             (@       �       �                    �?      �?             $@       �       �                    �K@���Q��?             @       �       �                    �H@�q�q�?             @        ������������������������       �                     �?        �       �                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     N@���Q��?             @       �       �                     M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?��l¿?�            �r@       �       �                   �U@�f��'�?�            �p@        ������������������������       �                     �?        �       �                    �R@�ߤ4u�?�            �p@       �       �                   �[@�Q����?�            �p@        �       �                   ph@�S����?             3@        ������������������������       �                     $@        �       �                    �K@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                    \@�w��c�?�            �n@        �       �                    �? 7���B�?5            @T@       �       �                    Z@0z�(>��?/            �Q@        ������������������������       �                     @@        �       �                   �k@$�q-�?            �C@        ������������������������       �                     5@        �       �                   �p@r�q��?             2@       �       �                    b@և���X�?             @       �       �                    �?      �?             @        ������������������������       �                      @        �       �                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     $@        �       �                    �D@@ o����?j            �d@        �       �                    b@r�q��?             @        ������������������������       �                     @        �       �                    �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @N@@��<W��?f            �c@       ������������������������       �        I            �\@        �       �                    �N@����?�?            �F@        �       �       	          `ff�?$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @@        ������������������������       �                      @        �       �                   @b@���!pc�?            �@@       �       �                    �?d}h���?             <@       �       �       	          ����?8�Z$���?             :@        �       �                   `]@���Q��?             @        ������������������������       �                      @        �       �                   0a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �^@���N8�?             5@        �       �                    @N@r�q��?             @        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                      @        �                          g@���Q��?             @       �                           �N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?              
                   �?�xGZ���?            �A@              	      
             �?���!pc�?             &@                                �?և���X�?             @                                �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                 `@�q�q�?             8@                                �Z@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @                    	          033�?��S���?	             .@        ������������������������       �                     @                                  M@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �t�b��
     h�h)h,K ��h.��R�(KMKK��hb�B0  �j�1N�?�J.g���?�)6���?6�����?W,<v���?S�����?�n���?~X�<��?;ڼOqɠ?\2�h��?              �?;�;��?;�;��?      �?                      �?�������?�������?�������?333333�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        ffffff�?333333�?      �?      �?      �?      �?              �?      �?              �?                      �?#
L:5�?r��+��?颋.���?]t�E]�?      �?      �?�������?xxxxxx�?              �?5�rO#,�?�{a���?      �?        l(�����?(������?�q�q�?9��8���?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?              �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        �������?�������?      �?      �?              �?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�m۶m��?%I�$I��?�m۶m��?�$I�$I�?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?���}�K�?��!XG�?��O��O�?l�l��?�$I�$I�?۶m۶m�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?        ���{��?�B!��?      �?              �?      �?۶m۶m�?�$I�$I�?      �?        /�袋.�?F]t�E�?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?        ��+2�?���\���?j�J�Z�?[�R�֯�?`��"���?����Mb�?ˠT�x�?���k��?      �?        UUUUUU�?UUUUUU�?�Mozӛ�?d!Y�B�?�q�q�?�q�q�?      �?      �?              �?      �?              �?              �?                      �?      �?      �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?GX�i���?���=��?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?        �?<<<<<<�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        z�rv��?~5&��?�?�������?�q�q�?�q�q�?              �?qG�w��?w�qGܱ?      �?        %I�$I��?۶m۶m�?              �?�Kh/��?h/�����?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?      �?        �������?�������?UUUUUU�?�������?�؉�؉�?ى�؉��?F]t�E�?/�袋.�?      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?              �?      �?                      �?      �?      �?�؉�؉�?ى�؉��?      �?      �?              �?      �?      �?              �?      �?                      �?l(�����?(������?              �?�������?�������?/�袋.�?F]t�E�?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?        ��A�:ܾ?H·�x$�?��[���?I����H�?�{a���?5�rO#,�?d!Y�B�?Nozӛ��?�?�������?�������?�������?              �?      �?      �?      �?                      �?�������?�������?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?              �?A�.��?x'Z���?~5&��?���¯�?      �?        3A�L-�?�4�.��?�E���?��=���?^Cy�5�?(������?              �?UUUUUU�?UUUUUU�?              �?      �?        �M!Д?Y��~Y�?h/�����?	�%����?H���@��?�ԓ�ۥ�?              �?;�;��?�؉�؉�?              �?UUUUUU�?�������?۶m۶m�?�$I�$I�?      �?      �?      �?              �?      �?      �?                      �?              �?              �?              �?�0�ӈ?�?�����?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ��N��y?�6b]z��?              �?l�l��?��I��I�?;�;��?�؉�؉�?      �?                      �?              �?      �?        t�E]t�?F]t�E�?۶m۶m�?I�$I�$�?;�;��?;�;��?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �a�a�?��y��y�?UUUUUU�?�������?      �?      �?              �?      �?                      �?              �?      �?        333333�?�������?      �?      �?      �?                      �?      �?        �A�A�?�_�_�?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?�q�q�?�q�q�?      �?                      �?�������?�?      �?        �q�q�?�q�q�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�c-hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK�h��B@<         �                    �?x��X���?C           ��@                                 �c@v��A���?4            ~@               
                   �`@�d����?U            @a@                                 �b@�K}��?;            �Y@       ������������������������       �        4            �V@               	       	          @33�?�C��2(�?             &@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                      
             �?�����H�?             B@       ������������������������       �                     7@                                   �?�	j*D�?
             *@                                  �?���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               }                   Pe@z����?�            `u@              :       	          pff�?{S"�?�            �t@               #       
             �?�s��:��?K            �\@                      	          833�?�+$�jP�?#             K@       ������������������������       �                     B@                                   @G@X�<ݚ�?             2@        ������������������������       �                     @                                   �?��S���?
             .@        ������������������������       �                     @                                  �_@���|���?             &@        ������������������������       �                      @               "                     O@�<ݚ�?             "@                                  �?���Q��?             @        ������������������������       �                      @                !                    �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        $       +                   `b@^n����?(             N@       %       *                    �? 	��p�?             =@        &       '                   �i@�q�q�?             @        ������������������������       �                      @        (       )                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     7@        ,       5                    �?`՟�G��?             ?@       -       0                   �]@8�A�0��?             6@        .       /                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        1       4                    �?$�q-�?	             *@        2       3                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        6       9                   �l@�����H�?             "@        7       8                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ;       l                   Xr@<J96���?�             k@       <       C                   `X@d#,����?l            �d@        =       >                   `W@���|���?             &@        ������������������������       �                     @        ?       B                    �?�q�q�?             @       @       A                   Pl@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        D       K                    �?XI�~�?d            @c@        E       J                   �`@�����H�?             2@        F       G       	             �?���Q��?             @        ������������������������       �                      @        H       I                   h@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        L       U                    j@�IєX�?Y             a@        M       T                    �?      �?             @@       N       O                   �\@PN��T'�?             ;@        ������������������������       �                     @        P       Q                   pb@ �q�q�?             8@       ������������������������       �                     5@        R       S                   g@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        V       c       	             @ ��WV�?A             Z@       W       X                   �m@F|/ߨ�?/            @T@        ������������������������       �                     =@        Y       \                   0n@ ��WV�?             J@        Z       [                    @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ]       b                    �?@�E�x�?            �H@       ^       _                   0c@��?^�k�?            �A@       ������������������������       �                    �@@        `       a                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        d       k       
             �?���}<S�?             7@       e       f                   8p@���7�?             6@       ������������������������       �                     *@        g       j                    �J@�����H�?             "@        h       i                     I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        m       n                   �r@      �?             J@        ������������������������       �                     @        o       t                    �?     ��?             H@        p       q                   �_@      �?              @        ������������������������       �                     @        r       s       
             �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        u       v       
             �?ףp=
�?             D@        ������������������������       �                     @        w       |                   @_@�?�|�?            �B@        x       {                   �t@z�G�z�?             @        y       z                    @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@        ~       �                    @K@���!pc�?	             &@              �                   �f@z�G�z�?             $@        �       �                   �b@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          `ff�?�	3��?           `{@       �       �       
             �?�L�x���?�            �s@        �       �                    �?��Q��?&             N@        �       �                    �?      �?
             (@       �       �                    T@ףp=
�?             $@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �b@      �?             H@       �       �                   �k@      �?             @@       �       �                   `X@ 7���B�?             ;@        �       �                   `Z@r�q��?             @       �       �                    V@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             5@        �       �                   c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          hff�?      �?
             0@       �       �                    �?X�<ݚ�?             "@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �G@؇���X�?             @        ������������������������       �                     @        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    X@�C͑V�?�            �o@        ������������������������       �                     �?        �       �                   0h@�U���?�            �o@       �       �                    �?0��kS֣?�            �o@       ������������������������       �        R             a@        �       �                    @M@@\�*��?D            @]@       �       �                   �]@�L��ȕ?4            @W@        �       �                   @d@@4և���?
             ,@        �       �                   �\@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        *            �S@        �       �                   ht@r�q��?             8@       �       �                   �c@�����?             5@       ������������������������       �        
             0@        �       �                   �]@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          ���@����v��?Q            �^@       �       �       
             �?b*0t��?C            �Y@       �       �                    �?` .�(�?1            �R@        �       �                   8p@���y4F�?             3@        ������������������������       �                     $@        �       �                    �?X�<ݚ�?             "@       �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�1�`jg�?&            �K@        �       �                   r@
;&����?             7@       �       �                    �?�t����?             1@       �       �       	          `ff�?d}h���?             ,@        ������������������������       �                     @        �       �                   �k@և���X�?             @        ������������������������       �                     @        �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?     ��?             @@       �       �                   P`@��<b���?             7@        �       �                   �b@����X�?             @       �       �                   �l@      �?             @        ������������������������       �                     �?        �       �                   `_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             0@        ������������������������       �                     "@        �       �                    �?\-��p�?             =@       ������������������������       �                     6@        �       �                   pb@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    `@R���Q�?             4@        ������������������������       �                     $@        �       �                    �?�z�G��?             $@       �       �                    l@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   0`@�q�q�?             @        ������������������������       �                     �?        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B  S��6�?ם,�d�?DDDDDD�?�������?)�3J���?��\;0��?�?�������?              �?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?�q�q�?              �?;�;��?vb'vb'�?�������?333333�?      �?                      �?              �?���?@���?�x��)�?<���u�?�k(���?��k(��?B{	�%��?/�����?              �?r�q��?�q�q�?      �?        �������?�?              �?]t�E]�?F]t�E�?              �?9��8���?�q�q�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?DDDDDD�?������?�{a���?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        �s�9��?�1�c��?颋.���?/�袋.�?�q�q�?�q�q�?      �?                      �?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?�h�?ڿ?�p	��?��[���?I����H�?F]t�E�?]t�E]�?              �?UUUUUU�?UUUUUU�?333333�?�������?      �?                      �?      �?        V~B����?5�wL��?�q�q�?�q�q�?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�?      �?      �?h/�����?&���^B�?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?;�;��?O��N���?�����H�?�Hx�5�?              �?;�;��?O��N���?UUUUUU�?UUUUUU�?      �?                      �?9/���?և���X�?�A�A�?_�_��?              �?      �?      �?              �?      �?                      �?d!Y�B�?ӛ���7�?F]t�E�?�.�袋�?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?      �?              �?      �?      �?      �?      �?        �������?333333�?              �?      �?        �������?�������?      �?        к����?*�Y7�"�?�������?�������?      �?      �?      �?                      �?              �?              �?F]t�E�?t�E]t�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?j�����?+���?;�S;�S�?+�+��?ffffff�?�������?      �?      �?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?      �?      �?      �?h/�����?	�%����?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?              �?      �?              �?      �?�q�q�?r�q��?�������?�������?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?�?�?              �?����|>�?��`0�?S��N^�?�5g"�<�?      �?        ���?^�^�?��~���?X`��?n۶m۶�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        �������?UUUUUU�?=��<���?�a�a�?      �?        333333�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?��/����?�h
���?�H%�e�?<�o�14�?��L���?�)�Y7��?6��P^C�?(������?      �?        r�q��?�q�q�?      �?      �?      �?                      �?              �?��)A��?��k߰�?�Mozӛ�?Y�B��?�������?�������?۶m۶m�?I�$I�$�?              �?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?��Moz��?��,d!�?�m۶m��?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?a����?�{a���?      �?        ۶m۶m�?�$I�$I�?              �?      �?        333333�?333333�?              �?333333�?ffffff�?�q�q�?9��8���?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$?mnhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM	hzh)h,K ��h.��R�(KM	��h��B@B         �                    �?TU�`��?P           ��@                                  `@Zw6G���?\           Ȁ@                                   @O@d۬����?<            @W@                                 0e@����p�?,             Q@                                  `@Hn�.P��?'             O@                     
             �?��(\���?             D@       ������������������������       �                     9@                                  �_@z�G�z�?	             .@       	                          @E@؇���X�?             ,@       
                           Z@$�q-�?             *@                                   @D@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@                                  �O@�q�q�?             @                                  \@z�G�z�?             @                                  `X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   �?�+e�X�?             9@                      	          ����?���Q��?             $@        ������������������������       �                      @                                  @L@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             .@                o       
             �?f�����?            �{@        !       T                    a@�ZbE���?^             a@       "       7                   �a@�W*��?A            @X@        #       (                   @\@��P���?            �D@        $       '                   �[@      �?              @       %       &                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        )       ,                    j@6YE�t�?            �@@        *       +                   h@      �?             @       ������������������������       �                     @        ������������������������       �                     @        -       .       	             �?�>����?             ;@        ������������������������       �                     *@        /       0       	          @33�?؇���X�?
             ,@        ������������������������       �                     �?        1       2                    �O@$�q-�?	             *@       ������������������������       �                     "@        3       6                   �s@      �?             @       4       5                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        8       9                   �b@���X�?$             L@        ������������������������       �                     $@        :       M                   p@�I� �?             G@       ;       B                   @_@�n`���?             ?@        <       =                    �?�IєX�?	             1@        ������������������������       �                     @        >       A                   �d@ףp=
�?             $@        ?       @       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        C       J                    �?X�Cc�?             ,@       D       E                   �b@�<ݚ�?             "@        ������������������������       �                     �?        F       G                   pe@      �?              @        ������������������������       �                     @        H       I                   �e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        K       L                   Pf@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        N       S       	          033�?���Q��?             .@       O       R                   xr@      �?	             (@       P       Q                    _@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        U       l       	          `ff@      �?             D@       V       e       	             �?�KM�]�?             C@        W       d                     R@z�G�z�?             .@       X       [                    �?؇���X�?             ,@        Y       Z                    `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        \       c                    �?�8��8��?
             (@       ]       ^       	          ����?؇���X�?             @       ������������������������       �                     @        _       `                    �?�q�q�?             @        ������������������������       �                     �?        a       b                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        f       g                    �?�nkK�?             7@       ������������������������       �        
             2@        h       i                   @_@z�G�z�?             @        ������������������������       �                      @        j       k       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        m       n                    @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        p       �                   �b@�yby��?�            0s@       q       �                    �?��O��"�?�            `q@        r       }                    �?"pc�
�?#            �K@        s       |                   f@�\��N��?             3@       t       {       	          ����?X�Cc�?
             ,@       u       v                   �^@�	j*D�?	             *@        ������������������������       �                     �?        w       x                   �_@      �?             (@       ������������������������       �                      @        y       z                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ~                          �s@������?             B@       ������������������������       �                     >@        �       �                    t@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @p����q�?�            �k@       �       �                    �? 9��?�            �j@       �       �                    �?�|���?l             f@        �       �                    �? �#�Ѵ�?            �E@       �       �                   �Y@������?            �D@        ������������������������       �                     �?        �       �                    ]@�(\����?             D@        �       �                   d@ףp=
�?             $@       �       �                    �H@      �?             @        ������������������������       �                      @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     >@        ������������������������       �                      @        ������������������������       �        S            �`@        ������������������������       �                    �B@        �       �                   �c@�z�G��?             $@       �       �                    �?؇���X�?             @       ������������������������       �                     @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   Pc@>���Rp�?             =@        �       �                     O@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���}<S�?             7@        ������������������������       �                      @        ������������������������       �                     5@        �       �                   @X@���_��?�            �w@        ������������������������       �                     @        �       �                    �?dlck+��?�            `w@       �       �       
             �?L������?�            s@       �       �                   P`@X��%�?�            Pp@        �       �                    �?���79��?B            @Y@       �       �                    �O@��|��?2            �S@       �       �       	          `ff�?ףp=
�?-            �Q@       �       �                    �?�������?             >@       �       �                    _@      �?             8@       ������������������������       �                     .@        �       �                   �_@�q�q�?             "@       �       �                   ``@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �K@�q�q�?             @       �       �                    �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     D@        �       �       	          ����?      �?              @        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        �       �                    �R@�(\����?g             d@       �       �                   �a@ � ���?e            �c@        �       �                    �?���7�?+            �P@        �       �                   �b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	             �?(;L]n�?%             N@        �       �                    @K@����X�?             @        ������������������������       �                     @        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        !            �J@        ������������������������       �        :             W@        �       �       	             @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@���!pc�?             F@       �       �                    �?д>��C�?             =@       �       �                    �?�d�����?             3@        ������������������������       �                     @        �       �                     K@�n_Y�K�?             *@        ������������������������       �                     @        �       �                   �^@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   �c@�q�q�?             @       �       �                    @N@z�G�z�?             @        ������������������������       �                      @        �       �                    \@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �       	             �?��S���?	             .@       �       �                    �N@�z�G��?             $@       ������������������������       �                     @        �       �                   �_@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@ٜSu��?.            @Q@       �       �                   Pj@��0{9�?            �G@        ������������������������       �                     9@        �       �                   �X@�X����?             6@        ������������������������       �                      @        �       �                    �?      �?             4@        ������������������������       �                      @        �       �                    �?r�q��?             2@       �       �                    q@      �?              @        ������������������������       �                     @        �       �       	          ����?���Q��?             @       �       �                    @M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �             
             �?�eP*L��?             6@       �       �                    @C@      �?             0@        ������������������������       �                     @        �                         0o@��
ц��?             *@       �                           L@      �?              @                                 �?���Q��?             @        ������������������������       �                      @                                �i@�q�q�?             @        ������������������������       �                     �?                    	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM	KK��hb�B�  ��Fc*�?y�\���?�p(���?	��*�?Hy�G�?7�p�7�?�����Ҳ?�������?�c�1ƨ?t�9�s�?333333�?�������?              �?�������?�������?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?      �?      �?              �?      �?                      �?      �?              �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?      �?        ���Q��?R���Q�?333333�?�������?              �?      �?      �?      �?                      �?              �?�5'��?���+c��?��髄��?16�='�?�Q�/�~�?_\����?�����?������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        e�M6�d�?'�l��&�?      �?      �?              �?      �?        h/�����?�Kh/��?              �?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?              �?      �?      �?      �?      �?      �?                      �?              �?۶m۶m�?I�$I�$�?      �?        Y�B���?Nozӛ��?�9�s��?�c�1��?�?�?      �?        �������?�������?�������?�������?              �?      �?              �?        %I�$I��?�m۶m��?9��8���?�q�q�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?              �?      �?        �������?333333�?      �?      �?      �?      �?              �?      �?              �?                      �?      �?      �?(�����?�k(���?�������?�������?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?        d!Y�B�?�Mozӛ�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�Q�}��?>r�dX�?i5	Q�E�?p�l�:��?/�袋.�?F]t�E�?y�5���?�5��P�?�m۶m��?%I�$I��?;�;��?vb'vb'�?      �?              �?      �?              �?      �?      �?      �?                      �?      �?              �?        �q�q�?�q�q�?      �?        �������?UUUUUU�?              �?      �?        C���RH�?������?��n��?��W[�:�?��.���?F]t�E�?�/����?�}A_Ч?p>�cp�?������?              �?333333�?�������?�������?�������?      �?      �?      �?              �?      �?      �?                      �?      �?              �?              �?              �?              �?        ffffff�?333333�?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �i��F�?GX�i���?UUUUUU�?�������?              �?      �?        ӛ���7�?d!Y�B�?              �?      �?        t�9G��?�Ƹ1n��?      �?        }�ٓ|�?�ʄm�?�Y�+���?�T�z�*�?��֡�l�? ��2)�?��g���?��N̓�?� � �?˷|˷|�?�������?�������?�������?�������?      �?      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?�������?�������?      �?                      �?              �?              �?�������?333333�?�&��jq�?ɞ��td�?F]t�E�?�.�袋�?UUUUUU�?�������?              �?      �?        �?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?      �?                      �?t�E]t�?F]t�E�?|a���?a���{�?y�5���?Cy�5��?              �?ى�؉��?;�;��?              �?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�?ffffff�?333333�?      �?              �?      �?              �?      �?                      �?%~F���?s��\;0�?L� &W�?m�w6�;�?              �?]t�E]�?�E]t��?      �?              �?      �?      �?        UUUUUU�?�������?      �?      �?              �?333333�?�������?      �?      �?              �?      �?                      �?              �?t�E]t�?]t�E�?      �?      �?              �?�؉�؉�?�;�;�?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��+hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@F         �       
             �?>���i��?R           ��@              u                   �b@��C���?F           X�@              h                    �?�L�j��?           �{@              %                    �?�=��=��?�            0s@                                   �?Np�����?!            �I@                      	          ���@�q�q�?             8@                                  �?��2(&�?             6@              	                    @E@d}h���?             ,@        ������������������������       �                      @        
              	          ����?�8��8��?             (@        ������������������������       �                     @                                  @q@      �?              @       ������������������������       �                     @                      	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                    �J@������?             ;@                                   �?�eP*L��?	             &@                                 `a@���Q��?             $@                                  �H@���Q��?             @        ������������������������       �                      @                                  Pn@�q�q�?             @        ������������������������       �                     �?                                  �s@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  `c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        !       "                    f@      �?             0@       ������������������������       �        	             ,@        #       $                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        &       [                   �a@     ��?�             p@       '       H                    �?4���|��?�             l@       (       9                    �? d���W�?n            @f@        )       0                    �?�:�^���?            �F@       *       +                   ``@Pa�	�?            �@@       ������������������������       �                     =@        ,       -       	             �?      �?             @        ������������������������       �                      @        .       /                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       6                    �K@      �?	             (@       2       5                    �?�����H�?             "@        3       4                   `Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        7       8                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        :       G                   �p@pJQg���?R            �`@       ;       @       	             �?XB���?:            �U@        <       =       	          ����?r�q��?
             (@       ������������������������       �                      @        >       ?                   �\@      �?             @        ������������������������       �                      @        ������������������������       �                      @        A       B                   �_@�}��L�?0            �R@       ������������������������       �        #            �L@        C       F                   g@�X�<ݺ?             2@        D       E                    b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     G@        I       L                   �T@��[�p�?            �G@        J       K                   �\@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        M       N                    i@�MI8d�?            �B@        ������������������������       �                     $@        O       R                    �?�<ݚ�?             ;@        P       Q                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        S       T                   �j@�LQ�1	�?             7@        ������������������������       �                      @        U       V                   �o@���N8�?             5@       ������������������������       �                     (@        W       Z                   �_@�����H�?             "@        X       Y                   �^@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        \       c                    �?r֛w���?             ?@        ]       b                    @      �?              @       ^       a                   @`@�q�q�?             @        _       `                    @L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        d       e                    �?�㙢�c�?             7@        ������������������������       �                     *@        f       g                   @Z@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        i       t       
             �?P#aE�?Q            �`@        j       o                   �a@�θ�?             :@       k       n       	          ����?�X�<ݺ?
             2@        l       m                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@        p       s       	          033@      �?              @       q       r                     O@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        B            �Z@        v       }                    �?�ҿf���?5            �T@        w       x       	          ����?     ��?             @@       ������������������������       �                     3@        y       z                    q@�θ�?	             *@       ������������������������       �                     "@        {       |                    b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ~       �                   pk@�\�u��?!            �I@               �                   �f@      �?             0@        �       �                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             (@        �       �                    @և���X�?            �A@       �       �                    �?J�8���?             =@       �       �                   �m@���!pc�?             6@        �       �                   �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             0@        �       �       	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?և���X�?             @       �       �                    �C@���Q��?             @        ������������������������       �                     �?        �       �                   e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	             �?r�q��?             @       �       �                    �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?z�G�z�?           �x@       �       �                    �?
��
�?�            �t@        �       �                    �?���Q��?A            �W@        �       �                    s@      �?             0@       ������������������������       �                     *@        �       �                    @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?bf@����?6            �S@       �       �                    `P@     ��?#             H@       �       �                   �]@p�v>��?"            �G@        �       �       	          ����?X�Cc�?             ,@       �       �                   �U@�q�q�?	             (@        ������������������������       �                     �?        �       �                   �[@���|���?             &@       �       �                    �?      �?              @        �       �                   g@z�G�z�?             @        ������������������������       �                     �?        �       �                   Pa@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �h@6YE�t�?            �@@        ������������������������       �        	             (@        �       �                   d@���N8�?             5@        ������������������������       �                     "@        �       �                   �^@�q�q�?	             (@        ������������������������       �                     @        �       �                    �?      �?              @        �       �                   f@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �`@���Q��?             @        ������������������������       �                     �?        �       �                   �d@      �?             @        ������������������������       �                     �?        �       �                   �e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �h@�4�����?             ?@        �       �                   �^@8�Z$���?             *@        ������������������������       �                     �?        �       �                   `_@�8��8��?             (@       ������������������������       �                     "@        �       �                   0a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @N@X�<ݚ�?             2@       �       �                    �?�q�q�?
             .@        �       �                    @I@      �?             @        ������������������������       �                      @        �       �                   �b@      �?             @       �       �                   @b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @K@�<ݚ�?             "@       ������������������������       �                     @        �       �                   �c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�7��?�            @m@        ������������������������       �        4            @S@        �                         �g@�e�B�?k            �c@       �       �                    �?��)�G��?j            �c@        �       �                    �?d}h���?             <@        �       �                   Pl@�C��2(�?             &@       ������������������������       �                     @        �       �                    �O@      �?             @       �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �d@�t����?             1@        ������������������������       �                     @        �       �                    q@؇���X�?             ,@       �       �       	          833@$�q-�?             *@       ������������������������       �        
             (@        ������������������������       �                     �?        ������������������������       �                     �?        �                           @     8�?V             `@       �       �                   @[@�â��,�?S             _@        �       �                    c@�8��8��?             (@        �       �                   0n@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �t@�h����?K             \@       �       �                    I@��wڝ�?I            @[@        �       �                    �J@؇���X�?             @        �       �       	          333�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        D            �Y@        �       �                   @`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                    	          ����?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                `c@�{r٣��?,            �P@                                V@�>$�*��?            �D@        ������������������������       �                     1@                                 �?      �?             8@       	      
                  @r@�IєX�?             1@       ������������������������       �        	             ,@                                 �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �`@����X�?             @        ������������������������       �                     @                                 �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                `R@�+e�X�?             9@        ������������������������       �                     @                                 �M@P���Q�?             4@       ������������������������       �                     2@                                 @O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  �Q��Q��?W�W��?���S@�?+�/�?� O	��?�7�}���?P�A�C�?��/��?PPPPPP�?______�?UUUUUU�?�������?��.���?t�E]t�?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?              �?      �?              �?      �?              �?                      �?{	�%���?B{	�%��?t�E]t�?]t�E�?333333�?�������?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?�������?      �?                      �?              �?      �?      �?              �?      �?      �?              �?      �?              �?     ��?�h$��W�?�r����?B�P�"�?�^��׽�?l�l��?}�'}�'�?|���?|���?              �?      �?      �?              �?      �?      �?              �?      �?              �?      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �qA��?s���7G�?�{a���?GX�i���?UUUUUU�?�������?              �?      �?      �?              �?      �?        O贁N�?�_,�Œ�?              �?�q�q�?��8��8�?�������?�������?              �?      �?                      �?              �?m�w6�;�?�
br1�?�������?333333�?              �?      �?        L�Ϻ��?��L���?              �?�q�q�?9��8���?      �?      �?      �?                      �?Y�B��?��Moz��?      �?        �a�a�?��y��y�?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?�B!��?���{��?      �?      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        d!Y�B�?�7��Mo�?              �?�������?333333�?      �?                      �?�qA��?�蛣o��?�؉�؉�?ى�؉��?�q�q�?��8��8�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�������?UUUUUU�?              �?      �?                      �?              �?Y1P�M�?S��rY�?      �?      �?              �?�؉�؉�?ى�؉��?              �?      �?      �?      �?                      �?�������?�?      �?      �?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?�rO#,��?|a���?F]t�E�?t�E]t�?UUUUUU�?�������?              �?      �?              �?      �?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?333333�?�������?              �?      �?      �?      �?                      �?              �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?6���#�?)sp�s�?333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?��&��j�?T:�g *�?      �?      �?ڨ�l�w�?L� &W�?�m۶m��?%I�$I��?�������?�������?      �?        F]t�E�?]t�E]�?      �?      �?�������?�������?              �?      �?      �?      �?                      �?      �?                      �?              �?'�l��&�?e�M6�d�?      �?        �a�a�?��y��y�?      �?        �������?�������?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?��RJ)��?���Zk��?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?r�q��?UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?9��8���?              �?�������?333333�?              �?      �?              �?        ��[��[�?�A�A�?      �?        ��� ܍�?A����?�[��[��?� � �?I�$I�$�?۶m۶m�?]t�E�?F]t�E�?      �?              �?      �?      �?      �?              �?      �?              �?        �������?�������?              �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?      �?                      �?              �?     ��?      �?:�s�9�?�c�1Ƙ?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?N��ش�?�,�M�ɂ?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?��|��?|���?�����?�18���?              �?      �?      �?�?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?        R���Q�?���Q��?              �?ffffff�?�������?      �?              �?      �?              �?      �?        �t�bub�OA     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��1hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�A         �                    �?�&���?R           ��@              Y       
             �?�9f��A�?`           ��@                      	          ����?����ث�?�            �k@                                   �?�����H�?3            @T@       ������������������������       �                     H@                                  �i@���!pc�?            �@@               
                    �?��
ц��?             *@               	                   p`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �H@�eP*L��?             &@        ������������������������       �                     @                                   �M@r�q��?             @                                   \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?ףp=
�?             4@                     
             �?"pc�
�?             &@        ������������������������       �                     �?                                  a@ףp=
�?             $@       ������������������������       �                     @                                  `a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@               0                    �?^�tD|��?[            �a@              /                   �a@�θ�?/            �S@                                  ]@�q�q�?              K@        ������������������������       �                     *@               "                    �?�>$�*��?            �D@                !       
             �?8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        #       $                   @^@      �?             <@        ������������������������       �                      @        %       .                   �`@���B���?             :@       &       -                    �?      �?             8@       '       ,                     P@z�G�z�?	             .@       (       +                    ]@$�q-�?             *@        )       *                    @I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     8@        1       X                   �e@     x�?,             P@       2       W                    �?~|z����?'            �J@       3       :                   pj@��C���?#            �G@        4       9       	          ���@"pc�
�?	             &@       5       8                   �f@ףp=
�?             $@        6       7                    @N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ;       @                    �?)O���?             B@        <       ?       	             �?      �?              @        =       >                   `X@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        A       R                   �c@և���X�?             <@       B       I                   �b@����X�?             5@        C       H       	          `ff�?      �?              @        D       E                     M@z�G�z�?             @        ������������������������       �                     �?        F       G                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        J       Q                    �K@8�Z$���?	             *@       K       L                   �^@���Q��?             @        ������������������������       �                      @        M       N                    �F@�q�q�?             @        ������������������������       �                     �?        O       P                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        S       T       	          833�?؇���X�?             @        ������������������������       �                     @        U       V                   pq@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        Z       ]                   `X@     ��?�             t@        [       \                   0d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ^       �       	             �?��XA%��?�            �s@       _       p                    �?�X�<ݺ?�            �p@        `       e                   d@���V��?             �F@       a       d       	          ����? 7���B�?             ;@       b       c                    �F@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �                     @        f       i                    �?�q�q�?             2@        g       h                   hq@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        j       o                   `b@d}h���?             ,@       k       n                   �i@�8��8��?
             (@        l       m                    �C@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        q       |                    @L@���
���?�             l@       r       u                   `R@����Oq�?u            �g@        s       t                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        v       w                   �k@ S5W�?r             g@       ������������������������       �        :            �V@        x       y                   �f@�eGk�T�?8            �W@       ������������������������       �        5             V@        z       {                   @b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        }       �       	          ����?r�q��?             B@       ~       �                   0d@؇���X�?            �A@              �                    b@�+$�jP�?             ;@       �       �                   �^@�8��8��?             8@        ������������������������       �                     @        �       �       	            �?�����H�?             2@       �       �       	          ����?��S�ۿ?             .@       �       �                   ps@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    `@֭��F?�?             �G@        �       �                    �?������?             .@        ������������������������       �                     "@        �       �                    g@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   Pb@     ��?             @@       �       �                   �a@����X�?             5@       �       �                    �?���y4F�?
             3@        ������������������������       �                     (@        �       �                    d@և���X�?             @       �       �                    @O@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    U@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�0&���?�            pw@        �       �       
             �?�zv�X�?             F@       �       �                    �J@4�2%ޑ�?            �A@        �       �                   �a@�q�q�?
             (@        �       �                    �?�q�q�?             @       �       �                    �I@���Q��?             @       �       �                    b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �]@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   hu@�nkK�?             7@       ������������������������       �                     2@        �       �                    �?z�G�z�?             @       �       �                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �       
             �?4c�O��?�            �t@       �       �                   �[@dkRk?�?�            pq@        �       �                    �?������?             >@       �       �       	          033@8�Z$���?             :@       �       �                   0i@H%u��?             9@       �       �                    �?�θ�?             *@        �       �       	             �?և���X�?             @        ������������������������       �                      @        �       �                   @`@���Q��?             @        ������������������������       �                      @        �       �       	             @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �R@h�U���?�             o@       �       �                   �b@/����?�            �n@       �       �                   �p@��<b�ƥ?�            �l@       �       �                   0p@��Q���?k            �d@       �       �                    �D@��惡�?f             d@        �       �                    �?      �?              @        �       �       	          ����?      �?             @       �       �                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   `f@`#`��k�?`             c@       �       �                    �?���=��?^            �b@       ������������������������       �        D            @]@        �       �                   �`@Pa�	�?            �@@       ������������������������       �                     8@        �       �                   pb@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        �       �                    �K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        -            �O@        �       �                    q@     ��?             0@       �       �                    _@ףp=
�?             $@        �       �                   c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �q@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �              	          ����?���3�E�?!             J@        �       �                   �`@�q�q�?             8@        �       �                   `c@�<ݚ�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �`@z�G�z�?
             .@        ������������������������       �                     @        �       �                     L@���!pc�?	             &@       ������������������������       �                     @        �       �                   �h@���Q��?             @       �       �                   �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                 �?h�����?             <@       ������������������������       �                     6@                                �`@r�q��?             @                                @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��hb�Bp  \�\��?R��Q���?�FV�a��?�rS�<��?�����?<��=v��?�q�q�?�q�q�?              �?t�E]t�?F]t�E�?�;�;�?�؉�؉�?      �?      �?      �?                      �?t�E]t�?]t�E�?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?�������?�������?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?      �?      �?                      �?              �?6���?�d�v�'�?�؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?�����?�18���?;�;��?;�;��?              �?      �?              �?      �?      �?        ى�؉��?��؉���?      �?      �?�������?�������?;�;��?�؉�؉�?      �?      �?      �?                      �?              �?      �?                      �?      �?                      �?     ��?      �?�	�[���?��sHM0�?L� &W�?g���Q��?/�袋.�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?9��8���?��8��8�?      �?      �?      �?      �?              �?      �?              �?        ۶m۶m�?�$I�$I�?�$I�$I�?�m۶m��?      �?      �?�������?�������?      �?              �?      �?              �?      �?                      �?;�;��?;�;��?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?              �?      �?             ��?      �?UUUUUU�?UUUUUU�?              �?      �?        �'�}4��?o�&\��?��8��8�?�q�q�?[�[��?�>�>��?	�%����?h/�����?�Mozӛ�?d!Y�B�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?2Tv����?߼�xV4�?��S�O��?�Zk��?      �?      �?              �?      �?        <����?@bw�#v?      �?        ��=�ĩ�?�X�0Ҏ�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?�������?UUUUUU�?۶m۶m�?�$I�$I�?/�����?B{	�%��?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?�������?�?�q�q�?�q�q�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?�F}g���?br1���?�?wwwwww�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?�m۶m��?�$I�$I�?6��P^C�?(������?      �?        ۶m۶m�?�$I�$I�?      �?      �?      �?                      �?              �?              �?]t�E�?F]t�E�?              �?      �?        �� �rh�?���S��?�袋.��?��.���?�A�A�?�������?�������?�������?UUUUUU�?UUUUUU�?�������?333333�?      �?      �?              �?      �?              �?                      �?�������?UUUUUU�?              �?      �?        d!Y�B�?�Mozӛ�?              �?�������?�������?      �?      �?              �?      �?                      �?      �?        ./ih�K�?�򒆶�?�Elo�?}Hw2��?�?wwwwww�?;�;��?;�;��?���Q��?)\���(�?�؉�؉�?ى�؉��?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?              �?        ��"NT��?�����?�M!Ф?��/����?d!Y�B�?��7��M�?\��l���?K��
�?V�	���?��/�Zg�?      �?      �?      �?      �?      �?      �?      �?                      �?              �?              �?p�pŊ?@�?��?O贁N{?�/��b��?              �?|���?|���?              �?�q�q�?�q�q�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?              �?      �?      �?�������?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        b'vb'v�?O��N���?�������?�������?�q�q�?9��8���?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?      �?        F]t�E�?t�E]t�?      �?        �������?333333�?      �?      �?      �?                      �?      �?        �$I�$I�?�m۶m��?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�+VahG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@=         n                    �K@�O(�.��?@           ��@              C                    �?�n�����??            @                     
             �?��x�E�?�            @v@                                   �?���ׁs�?8             Y@                                  q@��S�ۿ?	             .@       ������������������������       �                     ,@        ������������������������       �                     �?                      	          ����?�t����?/            @U@        	                           �E@@-�_ .�?            �B@        
                           �?8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                     8@                                  q@�q���?             H@                                  �?�99lMt�?            �C@        ������������������������       �                     @                      
             �?     ��?             @@                                   �?      �?              @                                 �\@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                      	          033�?�8��8��?             8@        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �                     "@               B       	          `ff @     p�?�             p@              3                    �?<��ٵ�?�            �o@               (                   i@P̏����?(            �L@               %                   �d@���Q��?             4@              $                    �?      �?
             ,@               !       	             �?�z�G��?             $@       ������������������������       �                     @        "       #                   `T@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        &       '                    �G@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        )       0                   �b@@-�_ .�?            �B@       *       +                   �b@Pa�	�?            �@@       ������������������������       �                     2@        ,       -                    �E@��S�ۿ?
             .@        ������������������������       �                     @        .       /                   @c@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        1       2                   po@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        4       ;                    �? %$��ݞ?w            �h@        5       :                   `e@      �?             @@       6       7                     H@�g�y��?             ?@        ������������������������       �                     0@        8       9                   �f@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        <       A                   @[@@�K�҈?g            �d@        =       @                   @c@�8��8��?             (@        >       ?                   �l@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        _             c@        ������������������������       �                     @        D       g                   �c@O�o9%�?f            �a@       E       H                   @Y@     |�?]             `@        F       G                   �[@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        I       f                    @��a�n`�?Y             _@       J       K                   @e@4Qi0���?X            �^@        ������������������������       �                    �C@        L       W                    �?H��?"�??             U@        M       V       	             �?      �?             (@       N       O                    �?�q�q�?             "@        ������������������������       �                      @        P       U                    �J@և���X�?             @       Q       T                   �a@�q�q�?             @       R       S                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        X       Y                   �e@�n���?4             R@        ������������������������       �                      @        Z       [                   �Z@hA� �?3            �Q@        ������������������������       �                     �?        \       e                    �?��.N"Ҭ?2            @Q@       ]       d                    �? ��ʻ��?1             Q@        ^       c                   �\@�X�<ݺ?             2@        _       b       	          ����?      �?             @       `       a                   `[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        ������������������������       �        $             I@        ������������������������       �                     �?        ������������������������       �                     �?        h       k                    �?d}h���?	             ,@        i       j                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        l       m                    �C@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        o       �                    �?�z�G��?           @z@        p       �       
             �?��.k���?,            @U@       q       �                    @P@�'N��?            �N@       r       }                    �?>a�����?            �I@        s       t                   @_@8����?
             7@        ������������������������       �                     @        u       |                    b@     ��?             0@       v       {                   �r@��
ц��?             *@       w       x       	             �?���Q��?             $@        ������������������������       �                     @        y       z                    @N@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ~       �                    �L@h�����?             <@               �                   �g@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             8@        �       �                   �c@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �       	          ����? �q�q�?             8@       �       �                     R@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        ������������������������       �                     "@        �       �       	          pff�?do@I�l�?�            �t@        �       �                   P`@���>4��?D             \@        �       �       	          833�?      �?"             J@       �       �       
             �?     ��?              H@       ������������������������       �                     @@        �       �                    �?     ��?             0@       �       �                   �]@"pc�
�?	             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��Q��?"             N@       �       �                    �?���Q��?            �F@       �       �                    �?     ��?             @@       �       �                     N@�����?             5@       �       �                    �?      �?	             0@        �       �                    �?      �?             @        �       �                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                    c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�eP*L��?             &@       �       �                   �p@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   `d@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        �       �       
             �?z�G�z�?	             .@        �       �                   �j@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �?�YK��?�            �k@       �       �                    c@�C��2(�?f            @c@       �       �                    �?�x�+���?`            @b@        �       �                    `@@�0�!��?             A@        �       �                   �^@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �P@H%u��?             9@       �       �                   @R@     ��?             0@        ������������������������       �                     �?        �       �       	          033@�r����?             .@       ������������������������       �        	             (@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �       
             �?���>4ֵ?J             \@       �       �                   pi@Pa�	�?A            �X@        �       �                    �?�����H�?             ;@       �       �                   `_@R���Q�?             4@       ������������������������       �                     .@        �       �       	             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        /             R@        �       �       	          033�?8�Z$���?	             *@       ������������������������       �                      @        �       �                   `b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    q@      �?              @       �       �                    �?r�q��?             @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �e@(���X�?+            @Q@       �       �                    _@j�'�=z�?)            �P@        �       �       
             �?      �?             (@        ������������������������       �                     @        �       �                   �a@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                   b@�{��?��?!             K@       �       �                   �b@(L���?            �E@       �       �                   �p@(;L]n�?             >@       ������������������������       �                     ;@        �       �                    �?�q�q�?             @       �       �                   Hr@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    d@�n_Y�K�?             *@        �       �                   �c@r�q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @N@�eP*L��?             &@        ������������������������       �                     @        �       �                   `c@r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �6S���?��rV��?T��cW�?W�ҋ8Q�?\���?ҏ~���?�(\����?��Q���?�������?�?      �?                      �?�������?�������?к����?S�n0E�?;�;��?;�;��?              �?      �?                      �?�������?�������?�o��o��?5H�4H��?      �?              �?      �?      �?      �?�������?333333�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?             ��?      �?�����?�SqК3�??���#�?��Gp�?�������?333333�?      �?      �?ffffff�?333333�?      �?              �?      �?              �?      �?                      �?UUUUUU�?�������?              �?      �?        S�n0E�?к����?|���?|���?      �?        �������?�?      �?              �?      �?              �?      �?              �?      �?              �?      �?        ������?և���X�?      �?      �?��{���?�B!��?      �?        �������?�?              �?      �?                      �?���|��?�����x?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?��RO�o�?�D+l$�?      �?     @�?      �?      �?              �?      �?        �c�1Ƹ?�s�9��?�On��?#6�a#�?              �?1�0��?�<��<��?      �?      �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?              �?              �?r�qǱ?r�q��?      �?        _�_�?���?      �?        ہ�v`��?�3J���?�?�������?�q�q�?��8��8�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?      �?              �?        I�$I�$�?۶m۶m�?      �?      �?      �?                      �?�������?�������?              �?      �?        333333�?ffffff�?�?�������?ާ�d��?�����?�?�������?8��Moz�?d!Y�B�?              �?      �?      �?�;�;�?�؉�؉�?�������?333333�?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?�������?�������?      �?                      �?�������?UUUUUU�?�������?�?      �?                      �?      �?        �bѲ
n�?�N�����?n۶m۶�?I�$I�$�?      �?      �?      �?      �?              �?      �?      �?/�袋.�?F]t�E�?      �?                      �?              �?      �?        �������?ffffff�?333333�?�������?      �?      �?=��<���?�a�a�?      �?      �?      �?      �?      �?      �?      �?                      �?      �?              �?        �������?�������?      �?                      �?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?;�;��?;�;��?              �?      �?        �������?�������?�������?333333�?              �?      �?              �?         �����?�����?F]t�E�?]t�E�?�4iҤI�?mٲe˖�?�������?ZZZZZZ�?UUUUUU�?UUUUUU�?              �?      �?        ���Q��?)\���(�?      �?      �?      �?        �?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�m۶mۦ?%I�$I��?|���?|���?�q�q�?�q�q�?333333�?333333�?              �?333333�?�������?              �?      �?                      �?              �?;�;��?;�;��?              �?�������?333333�?              �?      �?              �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        )�3J���?l�ځ��?|��|�?�|���?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        /�����?���^B{�?w�qG��?⎸#��?�?�������?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?ى�؉��?;�;��?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?]t�E�?t�E]t�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:�sdhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�G         �       
             �?������?9           ��@              +                    �?b��~T�?G           X�@                                   �c@V�K/��?2            �S@                                 �R@:���W�?(            �M@        ������������������������       �                     $@               	                   @[@և���X�?"            �H@                      	          ����?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        
              	          ����?      �?             D@                                   �?�C��2(�?             &@       ������������������������       �                     "@                                  �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                      	          ���@J�8���?             =@                                  `P@\X��t�?             7@                                 �n@�E��ӭ�?             2@        ������������������������       �                     @                                  �a@�q�q�?
             (@                                 �`@����X�?             @        ������������������������       �                     @                                  @b@      �?             @        ������������������������       �                     �?                                   �?�q�q�?             @                                  a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        !       "       
             �?z�G�z�?
             4@        ������������������������       �                     �?        #       *                    �?�S����?	             3@       $       %                   @_@�IєX�?             1@       ������������������������       �                     &@        &       )                   �o@r�q��?             @       '       (                    �I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ,       _                    �?��;D���?           �{@        -       <                    �?r֛w���?e            `c@       .       ;                    �?���!���?8            �S@       /       2       
             �?��k=.��?             �G@        0       1       	          ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       4       	          ����?:	��ʵ�?            �F@        ������������������������       �                     6@        5       8                   �^@�LQ�1	�?             7@        6       7                   �^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        9       :       	          ����?@�0�!��?             1@        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     @@        =       ^       	           33@��=A��?-             S@       >       C                    �?      �?,             R@        ?       B                    p@�q�q�?             2@       @       A                   �Z@؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     @        D       G                    @E@�E��ӭ�?$             K@        E       F       	          ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        H       [                   �c@��k=.��?            �G@       I       N                    �?,���i�?            �D@        J       M                    _@�θ�?	             *@        K       L       	          ���@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        O       Z                   �`@@4և���?             <@       P       Y                   @[@      �?
             0@       Q       X                    �N@"pc�
�?             &@       R       W                    �?ףp=
�?             $@       S       T                    �K@      �?              @        ������������������������       �                     @        U       V                   �^@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        \       ]                    �N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        `       �                   0c@t���:�?�            r@       a       �                    �?��(\���?�            �q@       b       �                    �?����˵�?�            �m@       c       l       	          ����?4����Y�?i            �e@        d       e       	          ����?4?,R��?             B@       ������������������������       �                     :@        f       g       	          hff�?      �?             $@        ������������������������       �                     @        h       k                    �?r�q��?             @       i       j                   �_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        m       �       	          033@PX�V|�?U            `a@       n                           �L@@\�*��?E            @]@       o       t                   `_@�[|x��?&            �O@        p       s                   �j@      �?             @@        q       r                   `Z@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     7@        u       x       
             �?��� ��?             ?@        v       w                    @H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        y       ~                    `@@4և���?             <@        z       }                   0j@���Q��?             @       {       |       	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     7@        ������������������������       �                     K@        �       �                   �Z@�C��2(�?             6@        ������������������������       �                     �?        �       �                   �\@���N8�?             5@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �        &            �N@        �       �       	          ����?�������?             F@        ������������������������       �                     *@        �       �       	          ����?¦	^_�?             ?@        �       �                     P@��S���?	             .@       �       �                    �J@�q�q�?             (@        �       �                    �H@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �N@؇���X�?             @        �       �                    b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@      �?             0@       ������������������������       �        	             ,@        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    _@X�<ݚ�?             "@        ������������������������       �                     @        �       �       	             @r�q��?             @       �       �                    q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �                           �?�Ҽݡ��?�            �x@       �       �                   @E@��,���?�            u@        �       �       	            �?      �?             @@        �       �                    �?��
ц��?             *@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?      �?              @       �       �                   `[@r�q��?             @        �       �                    @D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �       	          `ff�?�}�+r��?
             3@        �       �                    �?؇���X�?             @       �       �                   `a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �? *��X�?�            s@        �       �                    �? 1_#�?             �M@        �       �                    �?�q�q�?             8@        �       �                    d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �b@X�<ݚ�?	             2@        ������������������������       �                     @        �       �       	          @33�?�θ�?             *@       �       �                    @M@���!pc�?             &@       �       �                    @F@�����H�?             "@        ������������������������       �                     @        �       �                    �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                     L@(N:!���?            �A@       �       �       	          ����? �q�q�?             8@       �       �                    �?P���Q�?             4@        ������������������������       �                     @        �       �                   �d@��S�ۿ?	             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     @        �       �                     N@���!pc�?             &@        �       �                   `d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    @L@/����?�            �n@       �       �                    �?@�X��?�            `j@        �       �                   �b@���.�6�?             G@       �       �                    �?������?            �D@       �       �       	          ����?      �?             @@       �       �                   �_@���}<S�?             7@        �       �                   0c@r�q��?	             (@       ������������������������       �                      @        �       �                   d@      �?             @        ������������������������       �                     �?        �       �                   �d@�q�q�?             @        ������������������������       �                     �?        �       �                   0k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             &@        ������������������������       �                     "@        ������������������������       �                     "@        �       �                   �d@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        e            �d@        �       �                   p@z�G�z�?            �A@       �       �       	          ����? �q�q�?             8@       ������������������������       �                     4@        �       �                   �k@      �?             @       �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �P@�eP*L��?             &@       �       �                    �?      �?              @        ������������������������       �                     �?        �       �                   �`@؇���X�?             @        ������������������������       �                     @        �       �                   �p@      �?             @        ������������������������       �                      @        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �L@>n�T��?$             M@                                �B@�ʻ����?             A@        ������������������������       �                     @                                 �?���@M^�?             ?@                                @J@      �?             0@                               �e@8�Z$���?	             *@                               `b@�8��8��?             (@       ������������������������       �                     @        	      
                  �Z@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                    	             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     .@                    	          033�?r�q��?             8@                               0a@ףp=
�?             4@       ������������������������       �                     $@                                 �?z�G�z�?             $@                               �j@�����H�?             "@       ������������������������       �                     @                                �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                `U@      �?             @                                �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  �#@y��?'�_|C��?�Q�&���?�+U6S��?�Z܄��?�ґ=�?A�Iݗ��?_[4��?              �?۶m۶m�?�$I�$I�?�q�q�?�q�q�?      �?                      �?      �?      �?]t�E�?F]t�E�?      �?              �?      �?      �?                      �?|a���?�rO#,��?��Moz��?!Y�B�?r�q��?�q�q�?              �?�������?�������?�m۶m��?�$I�$I�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?      �?                      �?�������?�������?              �?(������?^Cy�5�?�?�?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�+c���?5'��P�?�B!��?���{��?T:�g *�?��	�Z�?br1���?g���Q��?      �?      �?      �?                      �?l�l��?��O��O�?              �?d!Y�B�?Nozӛ��?�������?UUUUUU�?              �?      �?        �������?ZZZZZZ�?      �?                      �?              �?������?(������?      �?      �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?              �?      �?                      �?r�q��?�q�q�?۶m۶m�?�$I�$I�?              �?      �?        br1���?g���Q��?8��18�?�����?�؉�؉�?ى�؉��?      �?      �?      �?                      �?              �?�$I�$I�?n۶m۶�?      �?      �?F]t�E�?/�袋.�?�������?�������?      �?      �?              �?�������?�������?      �?                      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        paRC4%�?ҳ�wY;�?333333�?�������?��/���?W'u_�?E'�危?�JC��?r�q��?�8��8��?              �?      �?      �?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?�&!��ȩ?��]tc�?^�^�?���?EQEQ�?]�u]�u�?      �?      �?�q�q�?�q�q�?      �?                      �?              �?�B!��?�{����?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?n۶m۶�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?F]t�E�?]t�E�?      �?        �a�a�?��y��y�?      �?      �?              �?      �?      �?      �?                      �?              �?              �?/�袋.�?t�E]t�?              �?�RJ)���?��Zk���?�?�������?�������?�������?�������?�������?              �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?�q�q�?r�q��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?e�����?�kNuA1�?Ğ���?���0��?      �?      �?�;�;�?�؉�؉�?�������?�������?      �?                      �?      �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        (�����?�5��P�?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?6����?R��ok��?	N�<�?��c+���?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?r�q��?      �?        �؉�؉�?ى�؉��?t�E]t�?F]t�E�?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?                      �?|�W|�W�?�A�A�?�������?UUUUUU�?ffffff�?�������?      �?        �������?�?      �?                      �?      �?        F]t�E�?t�E]t�?      �?      �?      �?                      �?      �?        ��/����?�M!Ф?��H����?�
��T�?���7���?Y�B��?p>�cp�?������?      �?      �?ӛ���7�?d!Y�B�?�������?UUUUUU�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?              �?        �������?�������?              �?      �?              �?        �������?�������?�������?UUUUUU�?      �?              �?      �?      �?      �?      �?                      �?      �?        ]t�E�?t�E]t�?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?      �?              �?      �?              �?        ��{a�?,�4�rO�?�������?<<<<<<�?              �?�s�9��?�c�1��?      �?      �?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?�������?�������?              �?�������?�������?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��hhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@D         �       	          ����?�lb���?@           ��@              9                    �?��c`��?/           �~@               (                    �?��}*_��?u            �g@              	       
             �?X3_��?Y            �a@                                   �? ,��-�?&            �M@                                   �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      J@        
       '                    �P@�0���?3            �T@              $                   �b@��مD�?1            @S@                                 �_@�㙢�c�?,            @Q@                                  �b@�4�����?             ?@                                  �?�}�+r��?             3@        ������������������������       �                     @                      	          ����?��S�ۿ?
             .@       ������������������������       �                     *@                                    N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?             (@        ������������������������       �                     �?                                   �?"pc�
�?             &@                                 @f@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?                                   �?�}�+r��?             C@                                  �r@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                #                    �?(;L]n�?             >@       !       "                    @N@���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        ������������������������       �                      @        %       &                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        )       0                   ``@��E�B��?            �G@       *       +       	          ����?(;L]n�?             >@       ������������������������       �                     :@        ,       -                    �E@      �?             @        ������������������������       �                      @        .       /                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        1       2                   Pj@�t����?
             1@        ������������������������       �                     "@        3       4                    �?      �?              @        ������������������������       �                     @        5       8       	          ����?���Q��?             @       6       7                   �t@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        :       o                    �?j��=k]�?�            �r@       ;       R                    @L@��B�5��?�            0p@       <       =                    �?��d5z�?�            `i@       ������������������������       �        E            �[@        >       K       
             �?��� ��?;            @W@        ?       J                    �?�5��?             ;@       @       A                    �?��H�}�?             9@        ������������������������       �                     $@        B       C                    �?���Q��?             .@        ������������������������       �                     @        D       I                   @`@      �?             (@       E       H                    �?      �?              @       F       G                   `]@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        L       M                    @G@����e��?.            �P@       ������������������������       �                    �F@        N       O                    m@���N8�?             5@       ������������������������       �        
             .@        P       Q                   �n@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        S       \       
             �?������?"             L@        T       Y                   `p@�E��ӭ�?             2@       U       X                   �_@؇���X�?	             ,@        V       W                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        Z       [       	          ����?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ]       j                   �b@�S����?             C@       ^       _                    �? 	��p�?             =@        ������������������������       �                     (@        `       g       	          ����?�t����?             1@        a       f                    �?r�q��?             @       b       c                   @c@      �?             @        ������������������������       �                      @        d       e                   p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        h       i                    �M@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        k       l                    ^@X�<ݚ�?             "@        ������������������������       �                     @        m       n                     P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        p       u                   �_@��Q��?             D@        q       r                    �?�z�G��?             $@        ������������������������       �                      @        s       t                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        v       y                    �G@�������?             >@        w       x                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        z       {       	          ���ٿ��2(&�?             6@        ������������������������       �                     �?        |       �                    �?�����?             5@        }       ~       
             �?z�G�z�?             $@        ������������������������       �                      @               �                   �`@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        �       �                    �?��Q��?           �z@        �       �                   pb@���g�?=            �Y@       �       �                    �O@�w��@�?#            �O@       �       �       
             �?���V��?            �F@       �       �                    @      �?             @@       ������������������������       �                     >@        ������������������������       �                      @        �       �                   �Y@�n_Y�K�?             *@        ������������������������       �                      @        �       �       	             �?���!pc�?             &@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?	             2@        �       �       
             �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          `ff�?z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �       	          033�?���Q��?             D@       �       �                    \@z�G�z�?             9@        ������������������������       �                      @        �       �                    �?�LQ�1	�?             7@        �       �                   0d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �e@P���Q�?             4@       ������������������������       �        
             3@        ������������������������       �                     �?        �       �                    �H@������?             .@        ������������������������       �                      @        �       �       	          033@8�Z$���?
             *@        �       �                   (p@���Q��?             @       �       �       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?6�����?�            pt@       �       �                   @f@@��ɨ�?�            �p@       �       �                    �?��c+��?�            �p@        �       �                   �`@�4�����?             ?@        �       �                    @N@��.k���?
             1@       �       �                   @_@�n_Y�K�?             *@        �       �                    @H@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?؇���X�?
             ,@        ������������������������       �                     �?        �       �                     K@$�q-�?	             *@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �Q@_k,D	�?�            �m@        ������������������������       �                      @        �       �       
             �?|�űN�?�            @m@        �       �       	          ����?�?�'�@�?             C@        ������������������������       �                     @        �       �                    �R@ >�֕�?            �A@       �       �                   �V@г�wY;�?             A@        ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                     �?        �       �                    @E@�ib�=�?�            �h@        �       �                   �b@�z�G��?	             $@       �       �                   �a@؇���X�?             @       ������������������������       �                     @        �       �                    �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	             �?�q�q�?             @       �       �                   �t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          ����?H��2�?x            @g@        �       �                    �?8��8���?             H@       �       �                    �?��� ��?             ?@       �       �                    @K@r�q��?             2@       ������������������������       �                     $@        �       �                   �_@      �?              @        ������������������������       �                     @        �       �                   �\@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �`@$�q-�?             *@        �       �                    �I@z�G�z�?             @        ������������������������       �                      @        �       �                    n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �k@�IєX�?	             1@       ������������������������       �                     &@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?��<b�ƥ?[            @a@       �       �                   0b@��V�I��?=            �W@       �       �       	          ����?`��>�ϗ?5            @U@        �       �                   @_@�X�<ݺ?             2@       ������������������������       �        	             ,@        �       �                     L@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        (            �P@        �       �                    �?�<ݚ�?             "@        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @M@؇���X�?             @       ������������������������       �                     @        �       �                   �n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     F@        ������������������������       �                     @        �                          �?��>4և�?#             L@       �                         `a@�G��l��?             E@        �                          @^@�8��8��?	             (@        ������������������������       �                     @                                 �F@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?d��0u��?             >@        ������������������������       �                     @                                 �?�+e�X�?             9@                   	          ���@��
ц��?             *@                                a@�eP*L��?             &@       	      
                   @I@X�<ݚ�?             "@        ������������������������       �                     @                                `^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �        
             ,@        �t�b��
     h�h)h,K ��h.��R�(KMKK��hb�B  �y�@$�?�4æ�m�?2�h�>�?��).��?B{	�%��?_B{	�%�?��V��?{2~�ԓ�?'u_[�?[4���?�$I�$I�?۶m۶m�?      �?                      �?              �?o4u~�!�?"�%��?��cj`��?�	qV~B�?�7��Mo�?d!Y�B�?���Zk��?��RJ)��?�5��P�?(�����?      �?        �������?�?      �?              �?      �?              �?      �?              �?      �?      �?        F]t�E�?/�袋.�?�������?�������?              �?      �?                      �?�5��P�?(�����?      �?      �?      �?                      �?�������?�?�.�袋�?F]t�E�?      �?                      �?      �?              �?      �?              �?      �?                      �?AL� &W�?�l�w6��?�?�������?              �?      �?      �?              �?      �?      �?              �?      �?        �������?�������?              �?      �?      �?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?)p�/�?\?"��C�?��i�}+�?A����?tl��?J��8D�?      �?        �{����?�B!��?h/�����?/�����?{�G�z�?
ףp=
�?      �?        �������?333333�?      �?              �?      �?      �?      �?      �?      �?              �?      �?                      �?              �?              �?�>����?|���?      �?        ��y��y�?�a�a�?      �?        �������?UUUUUU�?              �?      �?        I�$I�$�?n۶m۶�?r�q��?�q�q�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?                      �?(������?^Cy�5�?������?�{a���?      �?        <<<<<<�?�?�������?UUUUUU�?      �?      �?      �?              �?      �?      �?                      �?      �?        ]t�E�?F]t�E�?              �?      �?        r�q��?�q�q�?      �?        �������?�������?              �?      �?        �������?ffffff�?333333�?ffffff�?      �?              �?      �?      �?                      �?�������?�������?      �?      �?              �?      �?        ��.���?t�E]t�?              �?=��<���?�a�a�?�������?�������?      �?              �?      �?      �?                      �?      �?        ̳��<��?��0�?C����?^�	���?AA�?�}��}��?�>�>��?[�[��?      �?      �?              �?      �?        ى�؉��?;�;��?      �?        t�E]t�?F]t�E�?              �?      �?      �?      �?                      �?      �?      �?      �?      �?              �?      �?        �������?�������?      �?                      �?333333�?�������?�������?�������?              �?��Moz��?Y�B��?UUUUUU�?UUUUUU�?      �?                      �?ffffff�?�������?      �?                      �?�?wwwwww�?      �?        ;�;��?;�;��?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?4R1�:#�?s�3R1��?s�y�:�?�|�Э8�?��bk�غ?ʧ����?��RJ)��?���Zk��?�?�������?;�;��?ى�؉��?UUUUUU�?�������?              �?      �?              �?                      �?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?�������?�������?              �?      �?                      �?��c+���?����/��?      �?        ���?�������?y�5���?������?      �?        �A�A�?��+��+�?�?�?      �?                      �?      �?        /�����?����>4�?333333�?ffffff�?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        X`��?�~�駟�?�������?�������?�B!��?�{����?UUUUUU�?�������?              �?      �?      �?              �?333333�?�������?              �?      �?        ;�;��?�؉�؉�?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�?�?              �?UUUUUU�?�������?              �?      �?        d!Y�B�?��7��M�?AL� &W�?<�����?�?�������?�q�q�?��8��8�?              �?      �?      �?              �?      �?                      �?�q�q�?9��8���?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        I�$I�$�?۶m۶m�?1�0��?��y��y�?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?              �?      �?        wwwwww�?DDDDDD�?      �?        ���Q��?R���Q�?�؉�؉�?�;�;�?t�E]t�?]t�E�?�q�q�?r�q��?      �?        UUUUUU�?�������?      �?                      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJw�9hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         �                    �?�zܯ�V�?I           ��@              Q       
             �?��.��<�?^           �@                                   �?�>��+~�?�            �l@                                   �?��}*_��?!             K@                     	          ���@�7����?            �G@                                  b@RB)��.�?            �E@              
                    �?$G$n��?            �B@               	       	          ����?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@                                   �?PN��T'�?             ;@                                  �a@      �?             (@        ������������������������       �                     @                                  �_@���Q��?             @                                 @q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  `X@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@                      
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                      
             �? �ܽ��?j            �e@                      	          033@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @               N                    �Q@�1/z��?d            �d@               1                    �?B�xX�?b            `d@       !       ,                   pb@�IєX�?9            @U@       "       #                    �O@     ��?*             P@       ������������������������       �        !            �G@        $       +                   �`@�IєX�?	             1@       %       &                   @]@؇���X�?             @        ������������������������       �                     @        '       *                    �P@�q�q�?             @       (       )                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        -       .                    @L@��s����?             5@       ������������������������       �                     .@        /       0                   �c@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        2       M                   �s@����?)            �S@       3       L                   0o@�A+K&:�?(             S@       4       9                    �?Dc}h��?             L@        5       8       	          ����?      �?              @        6       7                   �_@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        :       E                   ``@r�qG�?             H@       ;       D                   `m@
j*D>�?             :@       <       C                    @O@�X����?             6@       =       B                    �?      �?             4@       >       A       	             @�q�q�?             (@       ?       @                   �k@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        F       K                     Q@�C��2(�?             6@       G       H                    @O@���N8�?             5@       ������������������������       �                     0@        I       J                   pk@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             4@        ������������������������       �                      @        O       P                    `R@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        R       �                    �?T�6|���?�            �s@       S       v                    @L@��.k���?�             q@       T       o                   �^@�X�<ݺ?�             k@        U       j       	            �?$�3c�s�?C            �W@       V       W                   �b@��p\�?:            �T@        ������������������������       �                     B@        X       c                    �?�LQ�1	�?"             G@        Y       ^                   d@      �?             $@        Z       ]                   �c@z�G�z�?             @       [       \                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        _       b                    ]@z�G�z�?             @       `       a                    e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        d       e                    �F@������?             B@       ������������������������       �                     7@        f       i                    o@$�q-�?	             *@        g       h                   @[@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        k       l                   �c@�q�q�?	             (@        ������������������������       �                     @        m       n                   �n@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        p       u                   �k@ ��7��?P            �^@        q       r                   �b@ �Jj�G�?"            �K@       ������������������������       �                    �I@        s       t                   �e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        .            �P@        w       �                   �c@���X�?$             L@       x       �                    @M@�㙢�c�?             G@        y       z                   @]@�n_Y�K�?	             *@        ������������������������       �                     @        {       |                   0b@X�<ݚ�?             "@        ������������������������       �                     @        }       ~                    �?�q�q�?             @        ������������������������       �                     �?               �       	          833@���Q��?             @       �       �                    �?      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @t@�C��2(�?            �@@       �       �                    �?      �?             @@        �       �                   �g@�<ݚ�?             "@        ������������������������       �                     @        �       �                   @d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     �?        �       �                    �?�z�G��?             $@        �       �                    �?؇���X�?             @       �       �       	          ����?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �O@�G�z��?             D@        ������������������������       �                     2@        ������������������������       �                     6@        �       �                   �b@:�ޟ���?�            �w@       �       �                    @�H�KY�?�            Pu@       �       �                    �?�.
�XX�?�            �t@        �       �                    �J@���#�İ?!            �M@        �       �       	             @�t����?
             1@       �       �                    a@      �?	             0@       ������������������������       �                     $@        �       �                   �a@r�q��?             @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     E@        �       �       	          ����? ���g=�?�            @q@       �       �                   �h@,�"���?l            @e@        �       �                   �_@@�j;��?4            �Q@       �       �       
             �?`Ql�R�?"            �G@       ������������������������       �                     C@        �       �       	             �?�����H�?             "@        �       �                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�q�q�?             8@       �       �                   pb@ףp=
�?             4@       ������������������������       �        
             .@        �       �       	             �?���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	             �?      �?             @       �       �                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Pi@�>�w��?8            �X@        ������������������������       �                      @        �       �       	             �?z�09JX�?7            @X@       �       �       
             �?�������?$             Q@       �       �       	          ����?�z�6�?             O@        ������������������������       �                     .@        �       �                    �?�7����?            �G@        �       �                    @I@r�q��?             (@        �       �                   �[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �\@">�֕�?            �A@        ������������������������       �                     @        �       �                   ``@z�G�z�?             >@        �       �                    �K@X�Cc�?             ,@        ������������������������       �                     @        �       �                    _@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	             �?      �?             0@        ������������������������       �                     �?        ������������������������       �                     .@        �       �                   �r@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     =@        �       �                    S@ �h�7W�?E            �Z@        �       �                    �J@�q�q�?             8@        �       �                   �Z@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?�KM�]�?             3@       ������������������������       �                     1@        ������������������������       �                      @        �       �                    �?����ȫ�?7            �T@       ������������������������       �        #            �K@        �       �                     K@ 7���B�?             ;@        �       �                    @J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     8@        �       �                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?�q�q�?             B@        �       �                    �H@�t����?             1@        �       �                   c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?�S����?             3@       �       �                    �?�t����?	             1@        �       �                   �q@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �f�f�?��L��L�?��W����?��P��|�?�r���?s���6��?_B{	�%�?B{	�%��?]AL� &�?G}g����?S֔5eM�?���)k��?к����?���L�?�������?�������?              �?      �?        &���^B�?h/�����?      �?      �?      �?        �������?333333�?      �?      �?      �?                      �?      �?        �������?�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�NV�#�?@l*9��?9��8���?�q�q�?      �?                      �?���\V�?��h���?��\w���?��(��I�?�?�?      �?     ��?              �?�?�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?�a�a�?z��y���?              �?UUUUUU�?UUUUUU�?      �?                      �?��-��-�?H�4H�4�?�k(���?y�5���?۶m۶m�?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?;�;��?b'vb'v�?]t�E]�?�E]t��?      �?      �?�������?�������?�m۶m��?�$I�$I�?      �?                      �?              �?              �?      �?              �?        F]t�E�?]t�E�?�a�a�?��y��y�?              �?�������?�������?              �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?'vb'vb�?b'vb'v�?�������?iiiiii�?��8��8�?�q�q�?1���\A�?x6�;��?�]�ڕ��?��+Q��?      �?        ��Moz��?Y�B��?      �?      �?�������?�������?      �?      �?              �?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        �q�q�?�q�q�?      �?        �؉�؉�?;�;��?�������?UUUUUU�?              �?      �?              �?        �������?�������?              �?      �?      �?      �?                      �?��:ڼ�?;ڼOqɀ?k߰�k�?��)A��?      �?              �?      �?      �?                      �?      �?        ۶m۶m�?I�$I�$�?�7��Mo�?d!Y�B�?;�;��?ى�؉��?      �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?        333333�?�������?      �?      �?      �?      �?              �?      �?              �?                      �?]t�E�?F]t�E�?      �?      �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?333333�?ffffff�?�$I�$I�?۶m۶m�?�������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?        �Z�&�?AiM~���?�r�!��?o���o�?䛌8j��?�l��?'u_[�?��N��?�?<<<<<<�?      �?      �?              �?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?                      �?ہ�v`��?��(�3J�?�������?�?H���@��?w�'�K�?W�+�ɕ?}g���Q�?              �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?UUUUUU�?�������?�������?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?      �?              �?      �?              �?        1ogH���?4$����?      �?        W?���?:*����?�������?�������?�Zk����?J)��RJ�?              �?G}g����?]AL� &�?UUUUUU�?�������?      �?      �?              �?      �?                      �?�A�A�?_�_��?      �?        �������?�������?�m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?              �?      �?              �?      �?      �?                      �?�������?UUUUUU�?      �?                      �?              �?"5�x+��?��sHM0�?�������?UUUUUU�?333333�?�������?      �?                      �?(�����?�k(���?              �?      �?        ������?������?              �?h/�����?	�%����?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�������?�������?�������?UUUUUU�?      �?                      �?              �?(������?^Cy�5�?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�whG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�?         `                   0`@x��X���?7           ��@                                  �d@�g�qT�?�            Pv@                                   �J@��b�h8�?O            �_@                                   �?��2(&�?             F@                                 @c@      �?             8@              	       
             �?��<b���?             7@                                   �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        
              
             �?R���Q�?             4@       ������������������������       �                     (@                      	             �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@                                   �M@ Df@��?3            �T@        ������������������������       �                     =@                                   @N@ 7���B�?             K@                                   [@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                  �]@���J��?            �I@       ������������������������       �                    �C@                                   �?�8��8��?             (@                                  �\@z�G�z�?             @        ������������������������       �                     @                      
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                C       	          pff�?��.۽0�?�            �l@        !       0                    �J@X�Cc�?4             U@        "       +                    �?�r����?             >@       #       *                    �?$�q-�?             :@        $       )                   pr@z�G�z�?             $@       %       (                   @\@�����H�?             "@        &       '                   �p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        ,       /                    �?      �?             @       -       .       
             �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        1       :                    �?|��?���?             K@        2       9                     R@     ��?             @@       3       8                    �?¦	^_�?             ?@       4       7                    ^@d}h���?             <@       5       6       
             �?�q�q�?	             2@        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     �?        ;       @       	          ����?���!pc�?             6@       <       =                   `q@�t����?             1@       ������������������������       �                     &@        >       ?                   �Z@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        A       B                   �^@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        D       I                    �?�F��O�?_            @b@        E       F                     L@      �?              @        ������������������������       �                     @        G       H                   `X@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        J       ]       
             �?p��%���?Y            @a@       K       L                   �e@���7�?V            �`@        ������������������������       �                     �?        M       R                    �?؀���˲?U            ``@        N       O                    �?�����?             5@       ������������������������       �                     2@        P       Q                    ^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        S       X       
             �?Ц�f*�?H            �[@        T       U                    �?      �?             0@       ������������������������       �                     $@        V       W                   @p@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        Y       \                   p`@��K2��?=            �W@        Z       [                    �?XB���?             =@       ������������������������       �                     <@        ������������������������       �                     �?        ������������������������       �        (            @P@        ^       _                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        a       �       
             �?���=�N�?U           ��@        b       �       	          ���@`џ�m�?�             m@       c       �                   �n@�8�jC��?k            `f@       d       �                    �?�Cc}��?D             \@       e       p                    �?�q���?8             X@        f       o                    �M@�ՙ/�?             E@       g       h                    �?�g�y��?             ?@        ������������������������       �                     $@        i       n                    �?����X�?             5@       j       k       
             �?�q�q�?             2@        ������������������������       �                     @        l       m                    �K@z�G�z�?             .@       ������������������������       �        	             (@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        q       �                   �c@��}*_��?             K@       r       s                    �?�+��<��?            �E@        ������������������������       �                     $@        t       {       	            �?4���C�?            �@@        u       z                   �l@r�q��?             (@       v       y                    �?�C��2(�?             &@        w       x                   pb@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        |       �                   �b@և���X�?             5@       }       ~                    I@      �?	             0@        ������������������������       �                     �?               �                    �?z�G�z�?             .@       �       �                   �`@���!pc�?             &@       �       �                   pb@�����H�?             "@        ������������������������       �                     @        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?�C��2(�?	             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   `a@     ��?             0@        ������������������������       �                     @        �       �                   �\@�z�G��?             $@        ������������������������       �                      @        �       �                    @M@      �?              @       ������������������������       �                     @        �       �                   @e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   Pb@h��Q(�?'            �P@        ������������������������       �                     ;@        �       �                    �?��Q��?             D@       �       �                    �?؀�:M�?            �B@       �       �                     P@|��?���?             ;@       �       �                    �L@���|���?             6@       �       �                    �G@�eP*L��?
             &@        ������������������������       �                     @        �       �                   �a@      �?              @       �       �                    �K@؇���X�?             @       ������������������������       �                     @        �       �                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     @        �       �                   @b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ���	@�>����?             K@       �       �                   `b@<���D�?            �@@       ������������������������       �                     1@        �       �                    �?      �?             0@       �       �                    �?؇���X�?             ,@        �       �       
             �?�q�q�?             @        ������������������������       �                      @        �       �                    c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             5@        �       �                    �?�i����?�            �t@       �       �                   @E@Tt�,b��?�            Pr@        �       �                    �?�ՙ/�?             5@        ������������������������       �                      @        ������������������������       �                     *@        �       �                   @g@������?�             q@       �       �                    �?�>����?�            �p@        �       �                    s@�x�E~�?8            @V@       ������������������������       �        -             R@        �       �                   s@�t����?             1@        ������������������������       �                     �?        �       �                   �d@      �?
             0@       ������������������������       �        	             .@        ������������������������       �                     �?        �       �       	          ����?����@��?u            �f@       �       �                    �?,�d�vK�?]            �a@        �       �                   �b@V������?            �B@       �       �                   �b@�'�`d�?            �@@        ������������������������       �        
             0@        �       �                    �?j���� �?             1@        �       �                     G@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    b@�z�G��?             $@       �       �                    �G@�<ݚ�?             "@       ������������������������       �                     @        �       �                   �c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        G            @Z@        �       �                    �?:�&���?            �C@        �       �                   �l@�q�q�?             (@        �       �                    �I@r�q��?             @        ������������������������       �                     @        �       �       	          hff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �c@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�>����?             ;@       �       �                   p@HP�s��?             9@       ������������������������       �        	             0@        �       �                   �p@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �       	          ����?�xGZ���?            �A@        �       �                    I@�t����?
             1@        ������������������������       �                      @        �       �                    �I@z�G�z�?	             .@        ������������������������       �                     "@        �       �                    �?      �?             @       �       �                   �c@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�<ݚ�?             2@       �       �                    �D@�	j*D�?             *@        ������������������������       �                      @        �       �       	          033�?"pc�
�?             &@       ������������������������       �                     @        �       �                   �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  S��6�?ם,�d�??�?��?9�]9�]�?�@ �?������?t�E]t�?��.���?      �?      �?��Moz��?��,d!�?UUUUUU�?UUUUUU�?              �?      �?        333333�?333333�?              �?      �?      �?      �?                      �?      �?                      �?��k���?c��7�:�?              �?h/�����?	�%����?UUUUUU�?UUUUUU�?              �?      �?        �?______�?              �?UUUUUU�?UUUUUU�?�������?�������?              �?      �?      �?      �?                      �?              �?&��~]�?m5x�@��?%I�$I��?�m۶m��?�������?�?�؉�؉�?;�;��?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?              �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        {	�%���?	�%����?      �?      �?��Zk���?�RJ)���?I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?              �?t�E]t�?F]t�E�?�?<<<<<<�?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?                      �?�P�B�
�?�իW�^�?      �?      �?              �?�������?�������?              �?      �?        ہ�v`��?�g��%�?F]t�E�?�.�袋�?      �?        �i��?h�T��?�a�a�?=��<���?              �?UUUUUU�?UUUUUU�?      �?                      �?�־a�?!O	� �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        W�+�Ʌ?��Q�٨�?�{a���?GX�i���?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��
hܭ�?��/G��?e�����?�����?�?d^J���?���}��?�$I�$I�?�m۶m��?�������?�������?�a�a�?�<��<��?�B!��?��{���?      �?        �$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?                      �?              �?_B{	�%�?B{	�%��?w�qG��?w�qG�?      �?        '�l��&�?m��&�l�?UUUUUU�?�������?F]t�E�?]t�E�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?�������?�������?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?]t�E�?F]t�E�?              �?      �?              �?      �?              �?333333�?ffffff�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        z�rv��?�Wc"=P�?              �?ffffff�?�������?v�)�Y7�?E>�S��?	�%����?{	�%���?F]t�E�?]t�E]�?t�E]t�?]t�E�?              �?      �?      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?/�袋.�?              �?      �?              �?        �������?�������?              �?      �?                      �?h/�����?�Kh/��?|���?|���?              �?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?                      �?��+Q��?�+Q��?��c�n-�?�*�L���?�a�a�?�<��<��?      �?                      �?iiiiii�?�������?�Kh/��?h/�����?����G�?p�\��?      �?        <<<<<<�?�?              �?      �?      �?      �?                      �?�C�rS��?��}kdu�?��9�h��?�z2~�Գ?�g�`�|�?o0E>��?6�d�M6�?'�l��&�?      �?        �������?ZZZZZZ�?۶m۶m�?�$I�$I�?              �?      �?        ffffff�?333333�?9��8���?�q�q�?      �?        333333�?�������?      �?                      �?              �?              �?      �?        �A�A�?�o��o��?�������?�������?�������?UUUUUU�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        �Kh/��?h/�����?q=
ףp�?{�G�z�?      �?        9��8���?�q�q�?              �?      �?              �?                      �?�A�A�?�_�_�?�������?�������?              �?�������?�������?      �?              �?      �?�������?333333�?      �?                      �?      �?        �q�q�?9��8���?;�;��?vb'vb'�?      �?        F]t�E�?/�袋.�?              �?      �?      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ@��hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�E         <                    �?�O(�.��?A           ��@               -       
             �?���N8�?x            �g@                                   @G@�l�]�N�?/             Q@                                    B@8�Z$���?
             *@        ������������������������       �                     �?                      	          ���@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        	       
                   �X@��N`.�?%            �K@        ������������������������       �                      @                                  �^@�q����?$            �J@                                   �J@X�<ݚ�?             "@        ������������������������       �                     @                                   �P@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               ,                    �?      �?             F@              +                    �Q@�q�q�?            �@@                                  �?¦	^_�?             ?@                                  �`@      �?              @        ������������������������       �                     @                                  @a@      �?             @        ������������������������       �                      @        ������������������������       �                      @               "                    �?8����?             7@              !                   u@z�G�z�?
             .@                                   �?$�q-�?	             *@                     	          ����?ףp=
�?             $@       ������������������������       �                     @                                   _@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        #       *       	             �?      �?              @       $       )                    @M@�q�q�?             @       %       (                   `b@z�G�z�?             @        &       '                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        .       7                    �?����&!�?I            @^@       /       6                    �?����q�?C            @[@        0       3                   �b@�����H�?             2@       1       2                   �s@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        4       5                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        7            �V@        8       9                   �`@�q�q�?             (@       ������������������������       �                     @        :       ;                   Hs@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =       �       
             �?��orf�?�           Ȇ@       >       }                   �a@R���Q�?           �{@       ?       z                    �R@h��jB�?�            0s@       @       Y                    �?�}�+r��?�             s@        A       F                    �?$�q-�?3            �S@        B       C                    �?      �?	             0@       ������������������������       �                     (@        D       E                   �]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        G       L       
             �?`Jj��?*             O@        H       K                    a@���Q��?             @       I       J                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        M       R                   `X@���U�?&            �L@        N       O                    �K@$�q-�?
             *@        ������������������������       �                      @        P       Q                   �W@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        S       T                   ``@`���i��?             F@       ������������������������       �                     =@        U       X                    �?��S�ۿ?             .@        V       W                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        Z       q                    ^@ \sF��?�            @l@       [       j       	          ����?ДXࣿ?W             a@        \       ]                   �i@�t����?+             Q@       ������������������������       �                     C@        ^       _       	          ����?������?             >@        ������������������������       �        	             ,@        `       a                    �J@      �?
             0@        ������������������������       �                     @        b       i                    �?���!pc�?             &@       c       h                     Q@z�G�z�?             $@       d       g                    �?�����H�?             "@       e       f                   �p@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        k       p                   @_@ ��ʻ��?,             Q@        l       m                   �^@P���Q�?             4@       ������������������������       �                     2@        n       o                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     H@        r       y                    �?�E�����?;            �V@       s       x                    \@P����?'            �M@        t       u                    �K@؇���X�?             @       ������������������������       �                     @        v       w       	          033�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        "             J@        ������������������������       �                     ?@        {       |                   pj@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ~       �                   �o@��}����?P            �`@              �                    �?|��?���?3            @T@        �       �                   �b@�+$�jP�?             ;@        �       �                   Pb@X�<ݚ�?             "@       �       �                   `X@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�X�<ݺ?             2@        �       �                   �`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �e@��}*_��?!             K@        �       �                   �d@�����H�?             "@       �       �                   `c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   ``@������?            �F@       �       �       	          ���@r�q��?             B@       �       �                    @��a�n`�?             ?@       �       �                   Pl@ȵHPS!�?             :@        ������������������������       �                     .@        �       �                   �\@���!pc�?             &@        ������������������������       �                     �?        �       �                    @J@z�G�z�?             $@        ������������������������       �                     @        �       �                   �b@�q�q�?             @        ������������������������       �                      @        �       �                    _@      �?             @       �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @_@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @O@�q�q�?             "@       ������������������������       �                     @        �       �                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   f@D>�Q�?             J@       �       �                    �?�:pΈ��?             I@        �       �       	          ���@��<b���?             7@       �       �       	          ����?؇���X�?             5@        �       �                    �I@�q�q�?             "@        ������������������������       �                     @        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        �       �                     M@�>����?             ;@       ������������������������       �        
             4@        �       �                    �?����X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	            �?��n���?�            r@       �       �                    �R@������?            `j@       �       �                    ]@4��?�?~             j@        �       �                   �b@�c�Α�?             =@       �       �                    �?��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        �       �                    �B@      �?	             ,@        ������������������������       �                     @        �       �                    �?���|���?             &@        �       �                    �E@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?D9���?k            `f@       �       �                    @L@8�Z� �?a            `d@       �       �                   �g@`o��b�?I             _@       ������������������������       �        H            �^@        ������������������������       �                     �?        �       �                   @c@8�Z$���?            �C@       �       �                   �c@ףp=
�?             >@       �       �                   @\@@4և���?             <@        �       �                   �^@�q�q�?             @        ������������������������       �                     @        �       �                   @`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     6@        �       �                   `n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     N@�q�q�?             "@       �       �                    c@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @E@     ��?
             0@        ������������������������       �                     �?        �       �                    h@������?	             .@        ������������������������       �                     @        �       �                    �I@�8��8��?             (@        ������������������������       �                     @        �       �                    @J@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �                          �?�{ /h��?3            �S@       �       �                    @E@z�J��?             �G@        ������������������������       �                     @        �                          �?�+��<��?            �E@       �       �       	          ����?�q�q�?             ;@        �       �       	          ����?r�q��?             (@        �       �                    ]@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �Z@��S���?             .@        �       �                   �]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�z�G��?             $@       �       �                    c@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �                           @K@      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?      �?             0@                    	          833�?z�G�z�?             @        ������������������������       �                     @                                �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              	                   @L@"pc�
�?             &@       ������������������������       �                     @        
                        @a@      �?             @        ������������������������       �                     �?                                �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 @L@�n`���?             ?@                                �X@�q�q�?             (@       ������������������������       �                     @        ������������������������       �                     @                                 �?�}�+r��?             3@       ������������������������       �        
             .@                                 �M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��hb�Bp  �6S���?��rV��?�a�a�?��y��y�?KKKKKK�?ZZZZZZ�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?                      �?� O	��?��oX���?      �?        �x+�R�?�Cj��V�?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?UUUUUU�?�RJ)���?��Zk���?      �?      �?              �?      �?      �?      �?                      �?8��Moz�?d!Y�B�?�������?�������?;�;��?�؉�؉�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?              �?      �?              �?              �?                      �?Sa���i�?���!pc�?���%�i�?�,�M�ɒ?�q�q�?�q�q�?�������?�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?�.sxQ��?�h�Cד�?333333�?333333�?|�x� �?hq���?(�����?�5��P�?;�;��?�؉�؉�?      �?      �?              �?      �?      �?      �?                      �?�B!��?���{��?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?p�}��?	�#����?;�;��?�؉�؉�?              �?�������?�������?              �?      �?        F]t�E�?F]t�E�?              �?�?�������?      �?      �?      �?                      �?              �?Vzja���?[X驅��?������?�������?�?<<<<<<�?              �?�?wwwwww�?              �?      �?      �?              �?F]t�E�?t�E]t�?�������?�������?�q�q�?�q�q�?�������?UUUUUU�?      �?                      �?      �?                      �?              �?�?�������?�������?ffffff�?              �?      �?      �?              �?      �?                      �?l�l��?P��O���?'u_[�?�V'u�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �qA��?8G�}s�?	�%����?{	�%���?B{	�%��?/�����?�q�q�?r�q��?�������?�������?      �?                      �?      �?      �?              �?      �?        �q�q�?��8��8�?UUUUUU�?�������?              �?      �?                      �?_B{	�%�?B{	�%��?�q�q�?�q�q�?      �?      �?              �?      �?                      �?wwwwww�?�?�������?UUUUUU�?�s�9��?�c�1Ƹ?��N��N�?�؉�؉�?      �?        F]t�E�?t�E]t�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �������?333333�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        vb'vb'�?b'vb'v�?�Q����?��Q���?��Moz��?��,d!�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?        h/�����?�Kh/��?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        RC4%�?��.k���?�.~��?w*���?�N��N��?ى�؉��?5�rO#,�?�{a���?�������?�?      �?                      �?      �?      �?              �?]t�E]�?F]t�E�?�������?�������?      �?                      �?      �?        Ų�����?�ir�y)�?���A2��?�Ŗ����?���{��?�B!��?      �?                      �?;�;��?;�;��?�������?�������?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?              �?      �?      �?              �?wwwwww�?�?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?                      �?�|˷|��?�A�A�?}g���Q�?AL� &W�?      �?        w�qG�?w�qG��?UUUUUU�?UUUUUU�?UUUUUU�?�������?�������?333333�?              �?      �?                      �?�������?�?�������?�������?              �?      �?        333333�?ffffff�?UUUUUU�?�������?              �?      �?              �?      �?      �?                      �?      �?      �?�������?�������?              �?      �?      �?              �?      �?        /�袋.�?F]t�E�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �c�1��?�9�s��?�������?�������?              �?      �?        (�����?�5��P�?              �?      �?      �?      �?                      �?�t�bub��;     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJث9hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@A         �                    �?��e�B��?E           ��@              =       	          ����?�Ee@���?7           �~@                      
             �?*L�9M�?s             f@                                  �b@H��?"�?7             U@                     	          ����?�#-���?/            �Q@       ������������������������       �        $            �K@                                   b@���Q��?             .@              	                    �?�q�q�?             "@        ������������������������       �                     @        
                          `^@���Q��?             @        ������������������������       �                     �?                                    L@      �?             @        ������������������������       �                     �?                                   `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                      	          ����?X�Cc�?             ,@                                 @c@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @                                   �?8����?<             W@                                  �d@�C��2(�?             6@                                  �?���N8�?             5@                                  �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        ������������������������       �                     �?               8                    �?<=�,S��?.            �Q@               %                   @E@�b��[��?#            �K@        !       $                     G@ףp=
�?             $@        "       #       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        &       +                    @F@�<ݚ�?            �F@        '       (                   �[@      �?             (@        ������������������������       �                     @        )       *                   pf@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ,       7                    @N@<���D�?            �@@       -       2                    �L@     ��?             @@       .       /                   `c@���7�?             6@       ������������������������       �                     4@        0       1                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       4                   �l@z�G�z�?             $@        ������������������������       �                     @        5       6                   p`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        9       <                   (p@��S���?             .@       :       ;                    b@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        >       y       
             �?tsrؚ��?�            �s@       ?       x                    �R@�E�J��?�            �p@       @       S                    �?���M�?�            �p@        A       H                   �_@     ��?             @@        B       G                    �?և���X�?             @       C       D                    �?      �?             @        ������������������������       �                     �?        E       F                   @[@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        I       P                   pc@H%u��?             9@       J       O                     K@���}<S�?             7@        K       N       	             �?      �?              @       L       M                   �p@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             .@        Q       R                    @O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                   �U@��!Dϸ?�            `m@        ������������������������       �                     @        V       Y                   �Q@���Rp�?�             m@        W       X                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Z       i                    ]@�94�s0�?�            �l@        [       ^                    �?<���D�?            �@@        \       ]                   �k@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        _       f                   �\@@4և���?             <@       `       e                    �? �q�q�?             8@        a       d                   �`@ףp=
�?             $@       b       c                   Pk@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     ,@        g       h                   `d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        j       w                   �i@��/�^�?z            �h@        k       n                   @X@F��}��?.            @R@        l       m                   �W@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        o       v                   pe@Pa�	�?)            �P@       p       q       	          033�?P���Q�?             D@       ������������������������       �                     :@        r       s       
             �?؇���X�?             ,@        ������������������������       �                     �?        t       u                    @G@$�q-�?             *@        ������������������������       �                     �?        ������������������������       �        
             (@        ������������������������       �                     :@        ������������������������       �        L             _@        ������������������������       �                      @        z       �                   �u@�%^�?            �E@       {       �                    �?z�G�z�?             D@        |       �                   �n@p�ݯ��?             3@       }       ~                    �?���|���?             &@        ������������������������       �                     �?               �                   �\@�z�G��?             $@        ������������������������       �                     �?        �       �                   �h@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �`@���Q��?             @        ������������������������       �                     �?        �       �                   0m@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �\@���N8�?             5@        �       �                    `@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                     @        �       �       
             �?n,
#9�?           �z@        �       �                    �?�'�7O��?j             e@       �       �                    �?�����?C            �Z@        �       �                    �?PN��T'�?             ;@       �       �                    �?HP�s��?             9@        �       �                   `n@      �?              @        �       �                    �?      �?             @       �       �                   �e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                      @        �       �                     Q@�2��?/            �S@       �       �                    �?p�}�ޤ�?,            @R@        �       �       	          ����?
j*D>�?             :@       �       �                   Pq@�q�q�?             5@       �       �                    �K@      �?             ,@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    ]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?t/*�?            �G@        �       �                    @I@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?��(\���?             D@        ������������������������       �                     @        �       �       	          ����?�8��8��?             B@       �       �                   @_@ȵHPS!�?             :@        �       �       	          ����?����X�?             @       �       �       	          ����?���Q��?             @       �       �                    �?      �?             @       �       �                    @J@�q�q�?             @        ������������������������       �                     �?        �       �                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�}�+r��?
             3@       ������������������������       �                     ,@        �       �       	          @33�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �e@r�q��?             @       �       �                    �R@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    \@d�;lr�?'            �O@        �       �                   p`@      �?              @       �       �                    �L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?X�;�^o�?"            �K@        �       �                     K@�θ�?             *@        �       �                   `c@      �?             @       �       �                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �`@�����?             E@       �       �                   �s@�g�y��?             ?@       ������������������������       �                     <@        �       �                   xt@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���!pc�?             &@       �       �                   �l@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    @L@�.^J��?�            Pp@       �       �                    I@�ʱ�O+�?z            �h@        �       �                    @���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�a�O�?v            @h@        �       �                   �d@�nkK�?             7@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �       �                   @[@ t�)Ї?g            `e@        �       �                    @G@      �?              @       ������������������������       �                     @        �       �                   `d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        a            `d@        �       �                    a@X��Oԣ�?*             O@        �       �                   `a@r�q��?             8@       ������������������������       �        
             .@        �       �                   @b@X�<ݚ�?             "@        ������������������������       �                      @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�˹�m��?             C@        ������������������������       �        
             2@        �                          @R���Q�?             4@       �                          b@      �?             0@       �       �                    �O@�����H�?             "@       ������������������������       �                     @        �                          �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                @`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�BP  �������?�������?q�����?�����?F]t�E�?]t�E]�?1�0��?�<��<��?_�_�?�A�A�?              �?�������?333333�?UUUUUU�?UUUUUU�?      �?        �������?333333�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?�m۶m��?%I�$I��?�������?�������?      �?                      �?      �?        d!Y�B�?8��Moz�?]t�E�?F]t�E�?��y��y�?�a�a�?      �?      �?      �?                      �?      �?                      �?�A�A�?X|�W|��?� O	��?־a��?�������?�������?      �?      �?      �?                      �?              �?9��8���?�q�q�?      �?      �?              �?      �?      �?      �?                      �?|���?|���?      �?      �?�.�袋�?F]t�E�?      �?              �?      �?      �?                      �?�������?�������?      �?              �?      �?              �?      �?                      �?�?�������?�q�q�?9��8���?              �?      �?              �?        ��o��o�?!� ��?��~���?�-���?�E(B�?��^����?      �?      �?۶m۶m�?�$I�$I�?      �?      �?              �?333333�?�������?              �?      �?                      �?���Q��?)\���(�?d!Y�B�?ӛ���7�?      �?      �?      �?      �?      �?                      �?              �?              �?      �?      �?      �?                      �?5���	%�?-�!c�]�?      �?        	�=��ܣ?O#,�4��?      �?      �?      �?                      �?���ϡ?��%���?|���?|���?�������?333333�?      �?                      �?�$I�$I�?n۶m۶�?UUUUUU�?�������?�������?�������?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?        n�%��ʔ?���;�Y�?����?��Ǐ?�?�$I�$I�?�m۶m��?              �?      �?        |���?|���?�������?ffffff�?              �?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?      �?                      �?              �?              �?      �?        �}A_�?�}A_��?�������?�������?Cy�5��?^Cy�5�?]t�E]�?F]t�E�?              �?ffffff�?333333�?              �?9��8���?�q�q�?      �?        333333�?�������?              �?      �?      �?              �?      �?                      �?�a�a�?��y��y�?      �?      �?              �?      �?                      �?      �?        !�n���?��"�{(�?��1G���?�g\��?\�琚`�?R�����?&���^B�?h/�����?q=
ףp�?{�G�z�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?                      �?�&��jq�?���JG�?�
*T��?�z��ի�?;�;��?b'vb'v�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�������?�������?              �?      �?        W�+���?�;����?�m۶m��?�$I�$I�?              �?      �?        333333�?�������?              �?UUUUUU�?UUUUUU�?�؉�؉�?��N��N�?�$I�$I�?�m۶m��?�������?333333�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?      �?                      �?(�����?�5��P�?              �?�������?�������?              �?      �?                      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        �eY�eY�?��i��i�?      �?      �?�������?�������?              �?      �?              �?        J��yJ�?�־a��?�؉�؉�?ى�؉��?      �?      �?      �?      �?      �?                      �?      �?                      �?�a�a�?=��<���?�B!��?��{���?              �?UUUUUU�?UUUUUU�?      �?                      �?t�E]t�?F]t�E�?�q�q�?�q�q�?      �?                      �?      �?        ��H���?��v��?}i�0V[�?gв�9��?333333�?�������?      �?                      �? tT����?����?�Mozӛ�?d!Y�B�?      �?      �?      �?                      �?      �?        ����?@��w?      �?      �?      �?              �?      �?              �?      �?              �?        c�1�c�?�s�9�?�������?UUUUUU�?      �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?              �?      �?        ��P^Cy�?^Cy�5�?      �?        333333�?333333�?      �?      �?�q�q�?�q�q�?      �?              �?      �?      �?                      �?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�E�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM	hzh)h,K ��h.��R�(KM	��h��B@B         �                   �b@X�<ݚ�?K           ��@              =                    �?�񴥑�?w           ��@               ,       
             �?$��r��?�            @o@               %                    �? d��0u�?N             ^@                                  �?b�2�tk�?0             R@                                  �u@؇���X�?             ,@                     	          pff�?$�q-�?
             *@        ������������������������       �                     @        	       
                   �Z@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   �K@�c�Α�?%             M@                                   g@д>��C�?             =@                      
             �?      �?              @        ������������������������       �                      @                      	             �?�q�q�?             @        ������������������������       �                      @                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                   �?���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@                                   @a@����"�?             =@                                 �\@���y4F�?             3@                                  �X@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @                                   �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        !       $                     N@�z�G��?             $@       "       #                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        &       +                    �?@��8��?             H@       '       *       	          ����?(;L]n�?             >@       (       )                   Hu@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     2@        -       6                   @c@z�G�z�?S            @`@        .       5                    @����e��?            �@@       /       4                    �P@f���M�?             ?@       0       3                    �?
j*D>�?             :@       1       2       	          ����?�G��l��?	             5@       ������������������������       �                     &@        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        7       8                    @M@�*v��?B            @X@       ������������������������       �        :             U@        9       <       	          hff�?��
ц��?             *@       :       ;                   �c@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        >       �                    @R@XT�z�q�?�            �s@       ?       P                   �[@|�`��?�            ps@        @       O                   �n@J�8���?             =@       A       J                    �?      �?             4@       B       I                   �i@�	j*D�?
             *@       C       H                   0a@"pc�
�?             &@       D       E                    ^@ףp=
�?             $@       ������������������������       �                     @        F       G                   @Y@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        K       L                    �?؇���X�?             @        ������������������������       �                     @        M       N       	          `ff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        Q       v       	          033�?heu+��?�            �q@       R       o       
             �?*~k���?b            �b@       S       T                   �i@t��ճC�?S            �`@        ������������������������       �        &             L@        U       f                    �?h�˹�?-             S@       V       W                   0j@��S�ۿ?$             N@        ������������������������       �                     �?        X       Y       	          hff�?����˵�?#            �M@        ������������������������       �                     2@        Z       a                   �[@��p\�?            �D@        [       \                   pm@r�q��?             (@        ������������������������       �                     �?        ]       `                   @_@�C��2(�?             &@        ^       _                   �t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        b       e                    @H@XB���?             =@        c       d                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     9@        g       n                    b@     ��?	             0@       h       i       	          ����?8�Z$���?             *@        ������������������������       �                     @        j       m       	          ����?�q�q�?             @        k       l                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        p       s       	          ����?�\��N��?             3@        q       r                     O@      �?              @       ������������������������       �                     @        ������������������������       �                     @        t       u                    �?���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        w       |                    �?�z�N��?[            ``@        x       {       	          033@$�q-�?	             *@       y       z                    �J@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        }       �                   �e@P����?R            �]@        ~       �       	             @�FVQ&�?            �@@              �                    �?���}<S�?             7@       �       �       
             �?�r����?             .@       �       �       	             �?$�q-�?
             *@        �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                    �E@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �        9            @U@        �       �                   �]@և���X�?             @       �       �                   �c@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?"f���r�?�            �u@        �       �                    �?$+ޠ�5�?C            @Z@       �       �                   �e@�f���?6            �T@       �       �                   ``@*O���?0             R@       �       �                    �?��s����?             E@        �       �                    �M@      �?              @       �       �                    �E@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   Xs@��hJ,�?             A@       �       �                    �E@<���D�?            �@@        �       �                     E@      �?             (@       �       �       
             �?ףp=
�?             $@       ������������������������       �                      @        �       �                    �C@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     O@���N8�?             5@       ������������������������       �        	             2@        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          `ff@���Q��?             >@       �       �                   d@�q�q�?             ;@       �       �                    �?     ��?             0@       ������������������������       �                     "@        �       �                    �?և���X�?             @        ������������������������       �                     �?        �       �                    c@      �?             @        ������������������������       �                      @        �       �                    �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�eP*L��?             &@        ������������������������       �                     @        �       �                    h@      �?              @        ������������������������       �                      @        �       �                    �M@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     6@        �             	             @.y����?�            �n@       �       �                    @L@h�˹�?�            �l@       �       �                   Ph@D9���?m            `f@       �       �                    �F@����!p�?k             f@        �       �                   �c@�Fǌ��?.            �S@        �       �                   `^@�}�+r��?             3@       �       �                    @E@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �        #             N@        �       �       	          ����?�$��y��?=            @X@       �       �                    �?Pa�	�?*            �P@       ������������������������       �        #             L@        �       �                    �?z�G�z�?             $@       ������������������������       �                     @        �       �       	          @33�?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    V@��a�n`�?             ?@        ������������������������       �                      @        �       �       	          ����?д>��C�?             =@        �       �                   �`@      �?             @       �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?HP�s��?             9@        ������������������������       �                     (@        �       �                     H@8�Z$���?	             *@        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�C��2(�?             &@       �       �                   @c@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �h@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          `ff�?~���L0�?            �H@       �       �                    @@�0�!��?             A@       �       �                    �L@�����H�?             ;@        �       �                   `f@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    c@�nkK�?             7@       ������������������������       �                     5@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                    �?���Q��?             @       �       �                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	             �?���Q��?             .@        ������������������������       �                     @        �       �                    �?�eP*L��?             &@        ������������������������       �                     @                                  �?      �?              @       ������������������������       �                     @        ������������������������       �                      @                                 `@@�0�!��?             1@        ������������������������       �                     "@                                 W@      �?              @        ������������������������       �                      @                    
             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM	KK��hb�B�  �q�q�?r�q��?$Zas ��?�RO�o��?�/�$�?�ʡE���?�������?DDDDDD�?9��8���?�8��8��?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?      �?        �������?UUUUUU�?              �?      �?                      �?�{a���?5�rO#,�?|a���?a���{�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�a�a�?��y��y�?      �?                      �?�i��F�?	�=����?(������?6��P^C�?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?        ffffff�?333333�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?�?�������?�?�������?              �?      �?                      �?              �?�������?�������?6�d�M6�?e�M6�d�?��Zk���?��RJ)��?;�;��?b'vb'v�?1�0��?��y��y�?      �?                      �?              �?              �?      �?        ���AG�? tT����?      �?        �;�;�?�؉�؉�?ffffff�?333333�?      �?                      �?              �?��c�^�?���3 ��?�E-����?AW o��?|a���?�rO#,��?      �?      �?;�;��?vb'vb'�?F]t�E�?/�袋.�?�������?�������?              �?      �?      �?              �?      �?              �?              �?        ۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?                      �?L� &W�?6�;���?�z=��?��^x/�?t�E]t�?�E]t��?              �?�5��P�?^Cy�5�?�?�������?      �?        ��/���?W'u_�?              �?��+Q��?�]�ڕ��?UUUUUU�?�������?      �?        F]t�E�?]t�E�?      �?      �?      �?                      �?              �?�{a���?GX�i���?      �?      �?      �?                      �?              �?      �?      �?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �5��P�?y�5���?      �?      �?      �?                      �?F]t�E�?]t�E]�?              �?      �?        ձ�6Ls�?qBJ�eD�?;�;��?�؉�؉�?UUUUUU�?�������?      �?                      �?              �?'u_[�?�V'u�?|���?>����?d!Y�B�?ӛ���7�?�?�������?;�;��?�؉�؉�?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?      �?                      �?              �?      �?      �?      �?                      �?              �?              �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        ������?��Tr��?�h��h��?�K��K��?�������?"�%��?�q�q�?�q�q�?�a�a�?z��y���?      �?      �?333333�?�������?              �?      �?                      �?�������?KKKKKK�?|���?|���?      �?      �?�������?�������?              �?      �?      �?      �?                      �?      �?        �a�a�?��y��y�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?      �?              �?      �?        ]t�E�?t�E]t�?              �?      �?      �?              �?�������?UUUUUU�?      �?                      �?              �?      �?                      �?v�[��?(2�ޟk�?^Cy�5�?�5��P�?Ų�����?�ir�y)�?/�袋.�?]t�E�?1���M��?�3���?�5��P�?(�����?�q�q�?�q�q�?      �?                      �?      �?              �?        ����?W?���?|���?|���?      �?        �������?�������?      �?        333333�?�������?              �?      �?        �c�1��?�s�9��?              �?a���{�?|a���?      �?      �?      �?      �?              �?      �?                      �?q=
ףp�?{�G�z�?      �?        ;�;��?;�;��?      �?      �?      �?                      �?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        ����>4�?������?ZZZZZZ�?�������?�q�q�?�q�q�?      �?      �?      �?                      �?�Mozӛ�?d!Y�B�?      �?              �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?333333�?              �?t�E]t�?]t�E�?              �?      �?      �?      �?                      �?�������?ZZZZZZ�?              �?      �?      �?      �?        UUUUUU�?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ!iTMhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�>         �       
             �?SH7�j�?J           ��@              -                    �?T��m�?J           ��@               (                   c@\��_��?1            �Q@                                  �?�eP*L��?(            �K@                     	          pff�?������?             ;@                                 �]@�q�q�?             5@                                   �?���Q��?             @        ������������������������       �                      @        	       
                   �R@�q�q�?             @        ������������������������       �                     �?                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?      �?             0@                     	          ����?������?
             .@        ������������������������       �                     @                                  �`@�q�q�?	             (@        ������������������������       �                      @                                   �I@z�G�z�?             $@                                   �?�q�q�?             @        ������������������������       �                     �?                                  �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                   �?�>4և��?             <@        ������������������������       �                     @                                   �H@���N8�?             5@        ������������������������       �                     @                '       	          ����?X�Cc�?	             ,@       !       &                    @      �?              @       "       %                   �`@����X�?             @        #       $                   0l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        )       ,       	          ����?     ��?	             0@        *       +                   �e@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        .       w                    �?�[s�&��?           �|@       /       l                   d@����Q8�?�            0v@       0       [       	          ����?p�_����?�             u@       1       V                    �?0G���ջ?{             j@       2       C                   `_@�7���?L             _@       3       8                    �?(�5�f��?0            �S@       4       5                    �O@����e��?'            �P@       ������������������������       �                     �K@        6       7                     P@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        9       :       
             �?8�Z$���?	             *@        ������������������������       �                     �?        ;       B       	          033�?�8��8��?             (@       <       =       	             �?r�q��?             @        ������������������������       �                      @        >       ?                   �Y@      �?             @        ������������������������       �                      @        @       A                   @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        D       O                    �?:	��ʵ�?            �F@       E       J                    `@4?,R��?             B@        F       G                    �E@���Q��?             $@        ������������������������       �                      @        H       I                     L@      �?              @       ������������������������       �                     @        ������������������������       �                      @        K       L                   �r@ ��WV�?             :@       ������������������������       �                     5@        M       N                   xt@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       U                    �?�q�q�?             "@       Q       R                    a@      �?             @        ������������������������       �                      @        S       T       	          ����?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        W       X                   Pz@ ��N8�?/             U@       ������������������������       �        ,             T@        Y       Z                   ``@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        \       ]                   �U@0�ޤ��?S            @`@        ������������������������       �                     �?        ^       _       	          033@ g�yB�?R             `@       ������������������������       �        =            �W@        `       a                    \@�IєX�?             A@        ������������������������       �                     �?        b       k                    �?Pa�	�?            �@@       c       d       
             �? ��WV�?             :@        ������������������������       �                     @        e       f                   8p@���N8�?             5@       ������������������������       �                     ,@        g       h                     J@؇���X�?             @       ������������������������       �                     @        i       j                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        m       t                   �`@�t����?             1@       n       o                   @d@d}h���?	             ,@        ������������������������       �                      @        p       q                     E@�8��8��?             (@        ������������������������       �                     @        r       s       	          ����?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        u       v                    �M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        x       �                    �?
io�v�?@            �Y@        y       z                    �K@�����?             C@        ������������������������       �                     (@        {       ~                   �`@��
ц��?             :@        |       }                     P@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@               �                   �l@     ��?
             0@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          033�?      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �B@�z����?+            @P@        �       �                   �f@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @Y@(��+�?(            �N@        �       �       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   pb@ܷ��?��?&             M@       �       �                   @^@`Ӹ����?            �F@        �       �                   �]@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �A@        �       �                   �q@�	j*D�?	             *@       �       �                    �?"pc�
�?             &@        ������������������������       �                     @        �       �                    _@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?@\�VK�?            Px@        �       �                    �?~31]���?X            @_@       �       �       	            �?�I{A�?F            �X@       �       �                    @O@���L��?1            �Q@       �       �                   �b@h��Q(�?.            �P@       ������������������������       �                    �B@        �       �                    �?��S���?             >@        �       �                   @d@      �?              @        �       �                    @L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �f@8�A�0��?             6@       �       �                    �?������?             1@       �       �                    ]@���|���?	             &@        ������������������������       �                     @        �       �                   �e@և���X�?             @       �       �                    �I@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?����"�?             =@        ������������������������       �                     @        �       �                    �J@�	j*D�?             :@        ������������������������       �                     @        �       �                    �?���Q��?             4@        �       �                    `@      �?              @        ������������������������       �                      @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @N@      �?	             (@        �       �                   �_@      �?             @        ������������������������       �                      @        �       �                   �a@      �?             @       �       �                   b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �a@ȵHPS!�?             :@       �       �                   ``@d}h���?
             ,@        ������������������������       �                     "@        �       �                    �I@���Q��?             @        ������������������������       �                      @        �       �                   h@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?�C��2(�?�            �p@        �       �                   @_@�|���?4             V@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                    [@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        0             T@        �       �                    �?D��2(�?t             f@       �       �                    c@�L���?d            �b@        �       �                    `@�q�q�?             2@        �       �                    �G@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                    c@P�2E��?]            @`@       �       �       	          pff�?���<_�?T            �]@       �       �                   @[@ pƵHP�?L             Z@        �       �                     H@      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �? �ׁsF�?H             Y@       �       �                    �O@�eGk�T�?E            �W@       ������������������������       �        B             W@        �       �       	          @33�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?@4և���?             ,@        �       �                   @e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    @      �?	             (@       �       �                   `c@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        �       �                   `R@��>4և�?             <@        ������������������������       �                     "@        �       �                   pp@�KM�]�?             3@       ������������������������       �                     1@        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ���t��?�~�E)�?��<b���?��p�F��?�K=��?$Zas �?t�E]t�?]t�E�?{	�%���?B{	�%��?UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?      �?�?wwwwww�?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?              �?�$I�$I�?�m۶m��?      �?        �a�a�?��y��y�?      �?        %I�$I��?�m۶m��?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?              �?      �?      �?      �?              �?      �?                      �?���!:ܿ?��λx�?��Vج?O�o�z2�?�θ�?ц�s��?�؉�؉�?vb'vb'�?��Zk���?)��RJ)�?�&��jq�?�=Q���?|���?�>����?              �?F]t�E�?]t�E�?      �?                      �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?      �?              �?      �?      �?              �?      �?                      �?l�l��?��O��O�?r�q��?�8��8��?�������?333333�?      �?              �?      �?              �?      �?        ;�;��?O��N���?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?                      �?�a�a�?�y��y��?              �?      �?      �?              �?      �?        z�z��?/�B/�B�?      �?        ����?�����?              �?�?�?      �?        |���?|���?;�;��?O��N���?              �?�a�a�?��y��y�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?�������?�������?۶m۶m�?I�$I�$�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?kch����?K��">��?Q^Cy��?^Cy�5�?      �?        �;�;�?�؉�؉�?�������?�������?              �?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?        �Z��Z��?[��Z���?      �?      �?              �?      �?        ;ڼOq��?q�����?UUUUUU�?UUUUUU�?      �?                      �?a���{�?��=���?l�l��??�>��?�������?�������?              �?      �?                      �?;�;��?vb'vb'�?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �N��&A�?�^�d��?���x�&�?V-��?[�R�֯�?K�Z�R��?��:��:�?_�_��?�Wc"=P�?z�rv��?      �?        �?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        /�袋.�?颋.���?�?xxxxxx�?F]t�E�?]t�E]�?              �?�$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?              �?      �?                      �?�i��F�?	�=����?      �?        ;�;��?vb'vb'�?              �?�������?333333�?      �?      �?              �?�������?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?              �?      �?      �?      �?              �?      �?                      �?              �?�؉�؉�?��N��N�?۶m۶m�?I�$I�$�?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?]t�E�?F]t�E�?��.���?F]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �E]t��?�袋.��?}���g�?L�Ϻ��?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?        _�^��?z�z��?+����/�?��/���?'vb'vb�?;�;��?      �?      �?      �?      �?      �?                      �?      �?        �G�z��?{�G�z�?��=�ĩ�?�X�0Ҏ�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?              �?      �?/�袋.�?F]t�E�?              �?      �?                      �?۶m۶m�?I�$I�$�?              �?�k(���?(�����?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ#EfghG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@D         |       	          ����?:���sQ�?=           ��@               c                    �?�r�k�h�?           �x@              6                    @L@�q����?�            @t@                     
             �?*��
�?�            @n@                      	          ����?�X����?$             F@                                  �?tk~X��?             B@               
                    �?�q�q�?             @              	                   �[@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  `X@ףp=
�?             >@                                  @`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                   �?`2U0*��?             9@       ������������������������       �                     2@                                    E@؇���X�?             @                                   �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                  �W@�X�<ݺ?�            �h@                                   �?�q�q�?             @                                  @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                -                    �?P�2E��?            `h@        !       *                    �?x�����?            �C@       "       )                   `\@؇���X�?            �A@        #       (                    �I@X�Cc�?	             ,@       $       '                    �?      �?             (@        %       &                    �G@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     5@        +       ,                   `\@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        .       /                    �?@f����?c            �c@       ������������������������       �        ;             Y@        0       5                   c@�h����?(             L@        1       4                   @[@`2U0*��?             9@        2       3                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     7@        ������������������������       �                     ?@        7       X                    �?D^��#��?8            �T@       8       ?                    �?�b��[��?$            �K@        9       :                    @M@��.k���?             1@        ������������������������       �                     @        ;       >                   �q@���!pc�?             &@       <       =                    @�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        @       C       
             �?�d�����?             C@        A       B       	          ����?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        D       E                   �Y@     ��?             @@        ������������������������       �                     �?        F       G                    �?��� ��?             ?@        ������������������������       �                     $@        H       I                    �L@��s����?             5@        ������������������������       �                      @        J       W                    �?�KM�]�?             3@       K       P                    �?�t����?             1@        L       O                    �O@z�G�z�?             @       M       N                   @g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Q       R                   pa@�8��8��?             (@        ������������������������       �                     @        S       T                    �N@z�G�z�?             @        ������������������������       �                      @        U       V                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        Y       b                   c@l��
I��?             ;@       Z       _                    @M@�ՙ/�?             5@        [       ^                   r@      �?              @       \       ]                   �^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        `       a       
             �?�θ�?
             *@       ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     @        d       y       	          833�?�1��u�?*            @R@       e       r                    �?�G�5��?&            @Q@       f       m                   �p@؇���X�?            �H@       g       l                   �d@��p\�?            �D@       h       i                   �a@P���Q�?             D@       ������������������������       �                     =@        j       k                   �b@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     �?        n       o                    �?      �?              @        ������������������������       �                      @        p       q                   �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        s       v                    �J@      �?             4@        t       u       
             �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        w       x                   �`@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        z       {                   `a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        }       �                   �b@�~���?5           H�@       ~       �       
             �?��Ç��?�            pz@              �                    �?��(�2Y�?�             w@        �       �                   �`@nM`����?             G@       �       �       	          ����?
j*D>�?             :@        ������������������������       �                     @        �       �                    �?D�n�3�?	             3@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�θ�?             *@        �       �                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @o@ףp=
�?             4@        �       �       	             �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        �       �                   0b@ wVX(6�?�            @t@       �       �                    �?��!�H�?�            Pr@        �       �       
             �?�חF�P�?"             O@        �       �                    �?�q�q�?             "@        ������������������������       �                     @        �       �                   �c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �H@�NW���?            �J@        �       �                   @_@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �O@@�E�x�?            �H@       ������������������������       �                     @@        �       �                   0k@�IєX�?             1@       ������������������������       �                     $@        �       �                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `P@P<��z4�?�            �l@       �       �       	          ����?�n����?y            �i@        �       �                   `j@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        �       �       	          033@@�~R(��?s            @h@       �       �                   �e@ ��N8�?d             e@       �       �                   @Y@��ϩ}��?a            �d@        �       �                    �?z�G�z�?             @       �       �                   Pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        ^             d@        �       �                   �g@�q�q�?             @       �       �                   @`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?ȵHPS!�?             :@        ������������������������       �                     @        �       �                   8p@R���Q�?             4@       ������������������������       �                     $@        �       �                   �\@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             8@        �       �                   �k@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �       	          033@r֛w���?             ?@       �       �                    �?�t����?             1@        �       �                     P@�q�q�?             @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �                   pb@և���X�?             ,@        ������������������������       �                     @        �       �       	          033@�eP*L��?             &@        ������������������������       �                     @        �       �                   @_@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @K@䯦s#�?#            �J@        �       �                    @I@X�<ݚ�?             ;@        �       �                    �?�θ�?             *@        ������������������������       �                      @        �       �                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?	             ,@       �       �                   `U@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    c@���B���?             :@       �       �                   �_@�LQ�1	�?             7@        ������������������������       �                     $@        �       �                   �`@�θ�?	             *@        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �c@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �                          �?f�Sc��?=            �X@       �       �       	             @��{�?6�?.            �R@       �       �                   r@�^����?%            �M@       �       �                   q@:�&���?            �C@       �       �                     M@l��\��?             A@       �       �                   �d@ 7���B�?             ;@       ������������������������       �        	             1@        �       �                    �?ףp=
�?             $@        �       �       	          033�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@����X�?             @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             4@        �                         �f@      �?	             0@       �             
             �?؇���X�?             ,@                                �`@      �?              @                               �\@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                    	          ����?��+7��?             7@        ������������������������       �                     �?        	                        �q@�GN�z�?             6@       
                         �?�t����?             1@        ������������������������       �                     @                                 q@�n_Y�K�?	             *@                                �F@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�b��B     h�h)h,K ��h.��R�(KMKK��hb�B  q���7T�?Ȏ �U�?V'�*6\�?T�᪓G�?ԭ�a�2�?�Hx�5�?�!pc��?�x?r���?]t�E]�?�E]t��?9��8���?r�q��?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?�������?�������?�������?333333�?      �?                      �?{�G�z�?���Q��?              �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?��8��8�?�q�q�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?_�^��?z�z��?��o��o�?�A�A�?۶m۶m�?�$I�$I�?%I�$I��?�m۶m��?      �?      �?�������?333333�?              �?      �?              �?                      �?      �?              �?      �?              �?      �?        �|˷|��?�A�Az?      �?        ۶m۶m�?�$I�$I�?���Q��?{�G�z�?      �?      �?              �?      �?              �?              �?        ,Q��+�?�]�ڕ��?� O	��?־a��?�?�������?              �?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?                      �?              �?Cy�5��?y�5���?UUUUUU�?�������?              �?      �?              �?      �?              �?�{����?�B!��?      �?        z��y���?�a�a�?              �?�k(���?(�����?<<<<<<�?�?�������?�������?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        h/�����?Lh/����?�a�a�?�<��<��?      �?      �?�������?UUUUUU�?              �?      �?                      �?�؉�؉�?ى�؉��?              �?      �?                      �?�1bĈ�?�s�Ν;�?�%~F��?��v`��?�$I�$I�?۶m۶m�?��+Q��?�]�ڕ��?�������?ffffff�?              �?F]t�E�?/�袋.�?      �?                      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�q�q�?�q�q�?              �?      �?        F]t�E�?/�袋.�?              �?      �?              �?      �?      �?                      �?d��ԗ3�?�Z�
3�?���E��?���.�?*�Y7�"�?�����?zӛ����?C���,�?b'vb'v�?;�;��?      �?        (������?l(�����?�������?UUUUUU�?      �?                      �?�؉�؉�?ى�؉��?      �?      �?      �?                      �?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�<ݚ�?k~X�<�?wury�?�|]����?��RJ)��?�Zk����?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �x+�R�?萚`���?      �?      �?      �?                      �?9/���?և���X�?              �?�?�?              �?�$I�$I�?۶m۶m�?              �?      �?        s�X�*�?yu�2^��?j6��bP�?�<����?;�;��?;�;��?              �?      �?        ���Id�?O"Ӱ�,�?�a�a�?�y��y��?�0��x?Ο��Y��?�������?�������?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�؉�؉�?��N��N�?              �?333333�?333333�?              �?333333�?ffffff�?      �?                      �?      �?      �?      �?      �?      �?                      �?              �?�B!��?���{��?�?<<<<<<�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?۶m۶m�?�$I�$I�?              �?t�E]t�?]t�E�?      �?              �?      �?      �?                      �?�V�9�&�?�����?r�q��?�q�q�?�؉�؉�?ى�؉��?              �?333333�?�������?              �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?ى�؉��?��؉���?Y�B��?��Moz��?              �?�؉�؉�?ى�؉��?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?����>�?������?�K~���?7�i�6�?u_[4�?W'u_�?�A�A�?�o��o��?------�?�������?	�%����?h/�����?      �?        �������?�������?      �?      �?              �?      �?              �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?              �?      �?              �?              �?      �?�$I�$I�?۶m۶m�?      �?      �?      �?      �?      �?                      �?              �?              �?      �?        Y�B��?zӛ����?      �?        ]t�E�?�袋.��?�������?�������?              �?ى�؉��?;�;��?�������?�������?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM	hzh)h,K ��h.��R�(KM	��h��B@B         �                   �b@�lb���?6           ��@                                 @E@䆎1�C�?�           ��@                                  �U@`Jj��?Z            `c@        ������������������������       �                     �?                      
             �?xJ��b,�?Y            @c@       ������������������������       �        F            �^@                                   �?¦	^_�?             ?@              	                    \@�ՙ/�?             5@        ������������������������       �                     @        
                           �?�E��ӭ�?             2@        ������������������������       �                     �?                                  �]@������?             1@        ������������������������       �                     @                                  @^@�q�q�?             (@                                   a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                                   �?؇���X�?             @                      	          hff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  �Z@ףp=
�?             $@                                  �X@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               -                    �F@�c�Q�?)           0~@               ,       
             �?:��?0            @V@               '                    �?���� �?            �D@              "                    `@�'�`d�?            �@@                !       	          `ff�?���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        #       &                   �Z@�LQ�1	�?             7@        $       %                    �C@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             3@        (       +                   �b@      �?              @       )       *                   0o@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     H@        .       w       
             �?n�ԉ	j�?�            �x@       /       n                    @4�S���?�            �p@       0       i                    �R@��FƘ��?�            �o@       1       X                   pn@����B��?�            �n@       2       ?                   �^@���-T��?N             _@        3       4                   �\@ 7���B�?#             K@        ������������������������       �                     �?        5       6                    �?�O4R���?"            �J@       ������������������������       �                     D@        7       8                    �?$�q-�?	             *@        ������������������������       �                     �?        9       >       	          ����?�8��8��?             (@        :       =                    �?z�G�z�?             @       ;       <                   `Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        @       A                   @Z@4�2%ޑ�?+            �Q@        ������������������������       �                      @        B       O                    �?H�V�e��?*             Q@       C       F                   �\@8��8���?             H@        D       E                   �a@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        G       L                    l@�7��?            �C@       H       K                    �?      �?             @@        I       J       	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        M       N                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       S                    @M@�G�z��?             4@       Q       R                    �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        T       W                   �`@�<ݚ�?             "@        U       V                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Y       Z                   �Q@ �q�q�?L             ^@        ������������������������       �                     �?        [       h                   �r@0x�!���?K            �]@       \       ]                   �Y@P���Q�?4             T@        ������������������������       �                     �?        ^       c                    �H@(�5�f��?3            �S@        _       `                   `@����X�?             @        ������������������������       �                     @        a       b       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        d       g       	            �?�k~X��?/             R@        e       f       	          ����?@4և���?             ,@       ������������������������       �                     *@        ������������������������       �                     �?        ������������������������       �        '             M@        ������������������������       �                    �C@        j       k       
             �?�<ݚ�?             "@        ������������������������       �                     @        l       m                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        o       v                   c@�q�q�?             (@       p       q                    �?      �?              @        ������������������������       �                     �?        r       s                   �[@����X�?             @        ������������������������       �                     �?        t       u       	          `ff @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        x       �       	          ����?<�I<���?S             `@       y       �                   �a@�*v��??            @X@       z       �                    `P@P��BNֱ?2            �T@       {       �                    �?�}��L�?.            �R@        |       �                    �?�8��8��?             (@       }       �                    �M@r�q��?             @        ~                          �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        (            �O@        �       �                    �P@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          ����?d}h���?             ,@       �       �                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        �       �       	          ����?     ��?             @@        �       �                   @b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?�eP*L��?             6@        �       �                     N@r�q��?             (@       ������������������������       �                     "@        �       �                    �?�q�q�?             @       �       �                   �n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @`@z�G�z�?             $@        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �p@��R[s�?�            �q@       �       �                   �O@>���a��?v            �f@        �       �                    �?�q�q�?             (@       �       �       	          ���
@���|���?             &@       �       �                    �?      �?              @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        �       �       	          `ff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `d@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �e@0,Tg��?n             e@       �       �       
             �?���O1��?m            �d@        �       �                    @G@��+7��?             G@        �       �                    �?�KM�]�?
             3@        ������������������������       �                      @        �       �                   Pf@"pc�
�?             &@       �       �       	          @33�?ףp=
�?             $@        �       �                    _@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ���@��}*_��?             ;@       �       �       	          ����?�q�q�?             8@        �       �                   �f@�q�q�?             @       �       �                   0e@z�G�z�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?r�q��?             2@       �       �       	          ����?�z�G��?             $@       �       �       	          hff�?      �?              @       �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   `]@ףp=
�?N             ^@        �       �                    �K@      �?             8@       �       �                   �Z@��<b���?             7@        ������������������������       �                     $@        �       �                    �G@�n_Y�K�?	             *@       �       �                    @E@X�<ݚ�?             "@       �       �                   pc@�q�q�?             @        ������������������������       �                      @        �       �                    f@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    l@      �?>             X@       �       �                    @M@\#r��?%            �N@       �       �                   �k@h�����?!             L@       ������������������������       �                    �J@        �       �                     G@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �A@        ������������������������       �                      @        �       �       
             �?Fx$(�?=             Y@        �       �                   Hr@�!���?             A@       �       �                    _@H%u��?             9@        ������������������������       �                     *@        �       �       
             �?      �?             (@        ������������������������       �                     �?        �       �                   pc@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �                          �L@�GN�z�?'            �P@       �                         @g@X�EQ]N�?            �E@       �                          �r@��p\�?            �D@        �       �                   �r@R���Q�?             4@       �       �                    �B@�KM�]�?             3@        �       �                     A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�IєX�?	             1@        �       �                    d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                      @                                 �?\X��t�?             7@                                 �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@                                r@      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KM	KK��hb�B�  �y�@$�?�4æ�m�?��9H��?�ےw�?�B!��?���{��?      �?        5�wL�?��8+?!�?              �?�RJ)���?��Zk���?�a�a�?�<��<��?      �?        r�q��?�q�q�?      �?        �?xxxxxx�?              �?UUUUUU�?UUUUUU�?333333�?�������?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?���C��?�
$޿�?S��Ԧ6�?Y�JV���?,Q��+�?jW�v%j�?'�l��&�?6�d�M6�?�������?333333�?      �?                      �?Y�B��?��Moz��?      �?      �?              �?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        @��DO��?`>�]X��?6��'��?z�6��?qК3[�?�ٝ4�?�y��!�?������?�RJ)���?[k���Z�?h/�����?	�%����?      �?        �x+�R�?:�&oe�?              �?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�A�A�?�������?      �?        ZZZZZZ�?iiiiii�?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?�A�A�?��[��[�?      �?      �?�������?�������?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?                      �?�������?�������?F]t�E�?/�袋.�?      �?                      �?9��8���?�q�q�?      �?      �?      �?                      �?      �?        UUUUUU�?�������?      �?        �5�5�?��~���?�������?ffffff�?      �?        �&��jq�?�=Q���?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?�q�q�?�8��8��?�$I�$I�?n۶m۶�?              �?      �?                      �?              �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?      �?              �?        sƜ1g��?4�9c��?���AG�? tT����?��FS���?���ˊ��?�_,�Œ�?O贁N�?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?              �?              �?      �?              �?      �?        I�$I�$�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�������?�������?              �?      �?        t�E]t�?]t�E�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�������?�������?      �?      �?              �?      �?                      �?X|�W|��?PuPu�?J��I���?؂-؂-�?UUUUUU�?UUUUUU�?F]t�E�?]t�E]�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?333333�?�������?      �?                      �?              �?              �?�0�0�?�<��<��?P�M�_�?���ˊ��?zӛ����?Y�B��?�k(���?(�����?      �?        /�袋.�?F]t�E�?�������?�������?      �?      �?              �?      �?              �?                      �?_B{	�%�?B{	�%��?�������?�������?UUUUUU�?UUUUUU�?�������?�������?      �?      �?      �?                      �?              �?      �?        �������?UUUUUU�?ffffff�?333333�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?�������?�������?      �?      �?��,d!�?��Moz��?      �?        ;�;��?ى�؉��?�q�q�?r�q��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?                      �?      �?      �?��:��?XG��).�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �������?�������?      �?                      �?      �?                      �?ףp=
��?R���Q�?�������?�������?���Q��?)\���(�?              �?      �?      �?      �?        F]t�E�?/�袋.�?      �?                      �?�q�q�?�q�q�?      �?                      �?�袋.��?]t�E�?w�qG�?qG�wĽ?�]�ڕ��?��+Q��?333333�?333333�?�k(���?(�����?      �?      �?      �?                      �?�?�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?                      �?!Y�B�?��Moz��?]t�E�?F]t�E�?              �?      �?              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJac�]hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK煔h��B�9         X       	          ����?��e�B��?F           ��@               #       
             �?�YE(\�?           �|@                                   �?��)�c{�?]             c@                                 �l@�nkK�?8             W@       ������������������������       �        &             Q@                                  �b@r�q��?             8@                                 xp@�}�+r��?             3@                                  �Z@ףp=
�?             $@        	       
                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@                                   c@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @               "                    �?��0u���?%             N@                                  �?�s��:��?             C@                      	          ����?r�q��?             (@                                  �?      �?              @                                  �J@؇���X�?             @       ������������������������       �                     @                                   �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   �?R�}e�.�?             :@        ������������������������       �                     @               !                   �^@�㙢�c�?             7@                                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     1@        ������������������������       �                     6@        $       ?                    �? ��om��?�            ps@        %       <                    �?d,���O�?:            �Y@       &       ;                    �P@z�G�z�?2            �V@       '       *                   �X@�T|n�q�?0            �U@        (       )                   �]@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        +       ,                   pc@�$�����?-            @T@       ������������������������       �                    �J@        -       .                    �?X�Cc�?             <@        ������������������������       �                      @        /       0                    @C@      �?             4@        ������������������������       �                      @        1       4                    �?X�<ݚ�?             2@        2       3                    ]@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        5       6                   �[@���!pc�?             &@        ������������������������       �                     �?        7       8                   �d@z�G�z�?             $@       ������������������������       �                     @        9       :                   �e@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        =       >                   @[@�q�q�?             (@        ������������������������       �                      @        ������������������������       �                     @        @       W                   �g@x�zKٲ?�             j@       A       L                    c@�ۛ�H@�?�            �i@       B       C                   pa@�1�:2�?w            @g@       ������������������������       �        W            �`@        D       K                   �a@ pƵHP�?              J@       E       J                    �?      �?             @@       F       I                   �c@ �q�q�?             8@        G       H                   @c@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �        	             ,@        ������������������������       �                      @        ������������������������       �                     4@        M       N                   Pc@z�G�z�?             4@        ������������������������       �                     �?        O       V                   �`@�S����?             3@        P       S                    �?և���X�?             @        Q       R                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        T       U                   p@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             (@        ������������������������       �                     @        Y       �       
             �?Ɲ��7P�?(           p|@       Z       u                    �?�������?�            �v@        [       t                   w@\�����?'            �K@       \       s                    �?r�q��?#             H@       ]       h                    �?�E��ӭ�?             B@       ^       _                   `X@R���Q�?             4@        ������������������������       �                     �?        `       g                    �?�KM�]�?             3@       a       b                   �]@z�G�z�?
             $@        ������������������������       �                     �?        c       d                   @q@�����H�?	             "@       ������������������������       �                     @        e       f                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        i       j                    �?     ��?             0@        ������������������������       �                     �?        k       r                   �s@��S���?
             .@       l       q                    �?�z�G��?             $@       m       n                   �`@�<ݚ�?             "@        ������������������������       �                     @        o       p       	          033�?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        v       �       	          ���@��|��?�            �s@       w       �                   �b@�P{6�I�?�             o@       x       �                    �?x��r��?�            `j@       y       |       	          ����?\���(�?a             d@        z       {                   p`@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @        }       �                    `R@ sAr�=�?\            �b@       ~       �                    �J@���g�X�?[            `b@               �                    @J@�*/�8V�?             �G@       �       �                    �?Du9iH��?            �E@       ������������������������       �                     B@        �       �                   �l@և���X�?             @        ������������������������       �                      @        �       �                    b@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?` A�c̭?;             Y@       �       �                    @L@�8���?"             M@        ������������������������       �                     :@        �       �                   pi@     ��?             @@        �       �                   @e@և���X�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     9@        ������������������������       �                     E@        ������������������������       �                     �?        �       �       	             �?��[�8��?             �I@        ������������������������       �                      @        �       �                    @M@Jm_!'1�?            �H@        ������������������������       �        
             1@        �       �       
             �?     ��?             @@        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    Y@������?             >@        ������������������������       �                      @        �       �                   �`@d}h���?             <@       �       �       	          ����?@4և���?
             ,@        �       �                   �p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �N@X�Cc�?             ,@        ������������������������       �                     @        �       �                   �[@"pc�
�?             &@        ������������������������       �                     �?        �       �                     P@ףp=
�?             $@        �       �       	          ����?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             C@       �       �                   �`@)O���?             B@       �       �                    X@$��m��?             :@        ������������������������       �                      @        �       �                    �H@�q�q�?             8@       �       �       	          ����?��S���?
             .@        ������������������������       �                      @        �       �                    �F@�n_Y�K�?	             *@       �       �                   x@���!pc�?             &@       �       �                   �o@�����H�?             "@       ������������������������       �                     @        �       �                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        �       �                   xr@z�G�z�?             $@       �       �       	          033�?�����H�?             "@        ������������������������       �                     @        �       �                   pc@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    j@ ������?(            �O@        �       �                   i@���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?        ������������������������       �                     E@        �       �                    ]@d�
��?>             V@        �       �                    �?�8��8��?	             (@        �       �                   pj@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �?��=A��?5             S@        �       �                    �?���"͏�?            �B@        ������������������������       �                     @        �       �                   `b@@�0�!��?             A@       ������������������������       �                     4@        �       �                   �s@և���X�?             ,@       �       �       	             �?���!pc�?             &@        ������������������������       �                     @        �       �                   �g@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ���@$�q-�?            �C@       �       �                    U@�}�+r��?             C@        ������������������������       �                     �?        �       �                    @�?�|�?            �B@       ������������������������       �                     ?@        �       �       	          033�?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �������?�������?�� њ��?���]���?��k(��?Cy�5��?d!Y�B�?�Mozӛ�?              �?UUUUUU�?�������?(�����?�5��P�?�������?�������?      �?      �?      �?                      �?              �?              �?333333�?�������?      �?                      �?""""""�?�������?�k(���?��k(��?�������?UUUUUU�?      �?      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �;�;�?'vb'vb�?      �?        d!Y�B�?�7��Mo�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�]i��?�����?�������?PPPPPP�?�������?�������?���)k��?6eMYS��?�������?�������?              �?      �?        uk~X��?X�<ݚ�?      �?        %I�$I��?�m۶m��?      �?              �?      �?      �?        �q�q�?r�q��?�m۶m��?�$I�$I�?              �?      �?        t�E]t�?F]t�E�?      �?        �������?�������?              �?�������?333333�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        
x>=n��?c,��?f�@*9�?C��ژ?�O?����?X`�v?      �?        'vb'vb�?;�;��?      �?      �?�������?UUUUUU�?�������?�������?      �?                      �?      �?              �?              �?        �������?�������?              �?(������?^Cy�5�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?      �?                      �?QQ�?x}�w}��?�ٸ�j�?�ɑA~��?A��)A�?߰�k��?UUUUUU�?UUUUUU�?�q�q�?r�q��?333333�?333333�?              �?�k(���?(�����?�������?�������?              �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?        �?�������?333333�?ffffff�?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?                      �?              �?� � �?˷|˷|�?����?�ҋ8Qy�?�
��T�?�^Fb5\�?�����̴?ffffff�?UUUUUU�?UUUUUU�?      �?                      �?*�Y7�"�?�`�|��?���+ݫ?��fG-B�?m�w6�;�?r1����?w�qGܱ?qG�w��?              �?۶m۶m�?�$I�$I�?              �?333333�?�������?      �?                      �?      �?      �?              �?      �?        ���Q��?
ףp=
�?a���{�?j��FX�?              �?      �?      �?۶m۶m�?�$I�$I�?�������?�������?      �?                      �?      �?                      �?              �?      �?        �������?�?      �?        ������?����X�?              �?      �?      �?      �?      �?              �?      �?        �?wwwwww�?      �?        ۶m۶m�?I�$I�$�?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?�m۶m��?%I�$I��?      �?        F]t�E�?/�袋.�?      �?        �������?�������?      �?      �?              �?      �?                      �?      �?      �?9��8���?��8��8�?�N��N��?vb'vb'�?              �?�������?�������?�?�������?              �?;�;��?ى�؉��?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �������?�������?�q�q�?�q�q�?              �?      �?      �?      �?                      �?      �?                      �?AA�?��}��}�?�a�a�?��y��y�?              �?      �?                      �?�袋.��?�.�袋�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?(������?������?*�Y7�"�?v�)�Y7�?      �?        �������?ZZZZZZ�?              �?۶m۶m�?�$I�$I�?t�E]t�?F]t�E�?              �?333333�?�������?              �?      �?              �?        �؉�؉�?;�;��?�5��P�?(�����?              �?*�Y7�"�?к����?      �?        �������?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJA�;6hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK텔h��B@;         �       
             �?Ly�'^��?C           ��@              '                    �?�s�?A           �@               &                   `d@�eP*L��?0            @S@                                  T@ꮃG��?,            @Q@        ������������������������       �                      @                                  �b@:2vz�M�?'            �N@                                  �?�J��%�?            �H@              	                    �?H%u��?             9@        ������������������������       �                     (@        
                           �?�θ�?
             *@                                  �?      �?              @                                 �m@����X�?             @       ������������������������       �                     @                                  0r@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  �b@r�q��?             8@                                 �l@�E��ӭ�?             2@                                  `a@���Q��?             @                                 �h@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                                   ]@8�Z$���?             *@                                    J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @                !                    f@r�q��?             (@       ������������������������       �                      @        "       %                    �?      �?             @       #       $       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        (       [                    �?8�Z$���?           �z@       )       D       	          ����?`-�I�w�?�             s@        *       +       	          833�?8��8���?W             b@       ������������������������       �        ,             Q@        ,       -                   �g@�=A�F�?+             S@        ������������������������       �                     @@        .       7                    @L@�X���?             F@        /       2                    �?�����H�?             2@        0       1                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        3       6                   p@      �?	             0@        4       5                   �m@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        8       =                   pm@      �?             :@        9       <                    i@�C��2(�?             &@        :       ;                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        >       C                    �?z�G�z�?             .@       ?       B                    �?�θ�?             *@       @       A       	            �?�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                      @        ������������������������       �                      @        E       Z                    �?      �?j             d@       F       K                   �Z@���tcH�?O            @^@        G       H       
             �?�q�q�?             @        ������������������������       �                     �?        I       J                    Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        L       O                   �e@���<_�?L            �]@        M       N                   @e@@-�_ .�?            �B@       ������������������������       �                    �A@        ������������������������       �                      @        P       Q                   Pa@ �)���?6            @T@        ������������������������       �                     B@        R       S                    @M@����?�?            �F@       ������������������������       �                     =@        T       U                   �p@      �?             0@        ������������������������       �                      @        V       W                    �?      �?              @        ������������������������       �                     @        X       Y                   �`@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                    �C@        \       �                   P`@������?P            @_@       ]       l                   �a@�Q����?1             T@        ^       i                     P@tk~X��?             B@       _       h                   �r@      �?             @@       `       c                    �?��a�n`�?             ?@        a       b                    �?      �?              @       ������������������������       �                     @        ������������������������       �                      @        d       e                    �K@�nkK�?             7@       ������������������������       �                     ,@        f       g                   `X@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        j       k       	          033@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        m       r                    W@v�X��?             F@        n       o                   �c@r�q��?             @       ������������������������       �                     @        p       q                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       |                   �o@���y4F�?             C@       t       u                   �l@ �Cc}�?             <@        ������������������������       �        	             (@        v       {                   �m@     ��?	             0@        w       z       	          `ff@      �?             @       x       y                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        }       �                   �p@      �?             $@       ~       �                   @_@z�G�z�?             @              �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �       	          `ff�?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?:	��ʵ�?            �F@        �       �                    �N@X�<ݚ�?             2@       �       �                    �J@      �?
             (@        �       �                   pb@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    p@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ;@        �       �       	            �?J��l��?           �y@       �       �                    I@X;h���?�            0s@        �       �                    �?
;&����?             7@        �       �                    �?�q�q�?             .@        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@       �       �                     P@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?����-��?�            �q@        �       �                    �?P�~D&�?,            �P@        �       �                     G@�G�z��?             4@        ������������������������       �                     @        �       �                    �?�	j*D�?
             *@       �       �                    �?؇���X�?             @       �       �                   �r@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @       �       �       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��0{9�?            �G@       �       �                    �I@(L���?            �E@       �       �                   �e@      �?             @@       ������������������������       �                     =@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    c@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        �       �                    @K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @L@�g�y��?�             k@       �       �                    �?�B:�g�?h            �e@       �       �                   �g@ A��� �?c            @d@       ������������������������       �        a             d@        �       �                    �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �                    �?(L���?            �E@        �       �                    @�q�q�?
             .@       �       �                   �`@r�q��?	             (@       ������������������������       �                     "@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pc@h�����?             <@       ������������������������       �        	             5@        �       �                   @`@؇���X�?             @        ������������������������       �                     @        �       �                   `q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �c@p�9�A��?H            @Z@        �       �       	          `ff�? >�֕�?            �A@        �       �                     O@      �?	             0@       ������������������������       �                     ,@        ������������������������       �                      @        ������������������������       �                     3@        �       �                    �?����X�?4            �Q@       �       �                   �`@�k�'7��?)            �L@       �       �       	          pff�?�z�G��?             >@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �L@�θ�?             :@       ������������������������       �                     3@        �       �                   �g@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �P@ 7���B�?             ;@       ������������������������       �                     9@        �       �                    @Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@�θ�?             *@        �       �                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ȫ�rV��?���T8�?�����?����֜�?]t�E�?t�E]t�?s��\;�?�%~F��?              �?��6�S\�?��!XG�?c}h���?9/����?)\���(�?���Q��?      �?        ى�؉��?�؉�؉�?      �?      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?r�q��?�q�q�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?�������?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?;�;��?;�;��?y�5�װ?Q^Cy��?�������?�������?              �?6��P^C�?��k(��?              �?�E]t��?]t�E�?�q�q�?�q�q�?      �?      �?              �?      �?              �?      �?UUUUUU�?�������?              �?      �?                      �?      �?      �?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?        �������?�������?�؉�؉�?ى�؉��?F]t�E�?]t�E�?      �?                      �?      �?                      �?      �?      �?�C��2(�?����|��?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        ��/���?+����/�?к����?S�n0E�?              �?      �?        �����H�?X�<ݚ�?              �?l�l��?��I��I�?              �?      �?      �?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?Zd;�O��?�MbX9�?ffffff�?�������?9��8���?r�q��?      �?      �?�c�1Ƹ?�s�9��?      �?      �?              �?      �?        d!Y�B�?�Mozӛ�?              �?�q�q�?�q�q�?      �?                      �?      �?              �?      �?      �?                      �?�.�袋�?颋.���?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?6��P^C�?(������?%I�$I��?۶m۶m�?      �?              �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?              �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?      �?                      �?l�l��?��O��O�?�q�q�?r�q��?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?UUUUUU�?      �?                      �?              �?>�Tr^�?��6���?��P�_?�?|�x� �?Y�B��?�Mozӛ�?UUUUUU�?UUUUUU�?              �?r�q��?�q�q�?�m۶m��?�$I�$I�?      �?                      �?              �?      �?      �?      �?                      �?ܥ���.�? �
���?kL�*g�?*g��1�?�������?�������?              �?vb'vb'�?;�;��?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?              �?      �?      �?      �?      �?                      �?              �?m�w6�;�?L� &W�?⎸#��?w�qG��?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?t�E]t�?]t�E�?      �?                      �?      �?      �?              �?      �?        ��{���?�B!��?��f���?Ȥx�L�w?,R�n��?�����Hy?      �?              �?      �?      �?                      �?      �?        ⎸#��?w�qG��?UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�m۶m��?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �? �����?p'p'�?�A�A�?��+��+�?      �?      �?              �?      �?                      �?�m۶m��?�$I�$I�?-����b�?Lg1��t�?ffffff�?333333�?      �?      �?      �?                      �?ى�؉��?�؉�؉�?      �?        �$I�$I�?۶m۶m�?      �?                      �?	�%����?h/�����?      �?              �?      �?              �?      �?        �؉�؉�?ى�؉��?      �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJkpkwhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�G         2                    �?x��X���?C           ��@               %       
             �?� !!��?w            �g@                                   �?��+��?2            �R@                                  �?x�����?            �C@                                 �b@(N:!���?            �A@        ������������������������       �        
             .@                      
             �?z�G�z�?             4@        ������������������������       �                     �?        	                          �c@�S����?             3@       
                           �N@և���X�?             @                                  �I@���Q��?             @        ������������������������       �                     �?                                   b@      �?             @                                  �K@�q�q�?             @        ������������������������       �                     �?                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     @                                  �g@؇���X�?            �A@                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?               "                   �u@     ��?             @@              !                   @m@��S�ۿ?             >@                                     K@"pc�
�?             &@                                 �j@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        
             3@        #       $                   @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        &       )                    T@ ���J��?E            @]@        '       (                   @b@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        *       1       	          ����?���͡?C            @\@       +       0                    �?�(\����?1             T@        ,       -                    s@؇���X�?
             ,@       ������������������������       �                     $@        .       /                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        '            �P@        ������������������������       �                    �@@        3       �                    �?���V��?�           ��@       4       _                    `@2��˕�?�            @y@        5       V                   c@*c̕6�?6            �U@       6       9                    �C@8�Z$���?0            �S@        7       8                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        :       Q       	             @      �?,             R@       ;       P                    �?��IF�E�?'            �P@        <       O                   �O@�q�q�?             8@       =       >       	          ������q�q�?             5@        ������������������������       �                      @        ?       H       	          ����?�d�����?             3@       @       G                    `@z�G�z�?             .@        A       F                    �?և���X�?             @       B       C                   `Y@���Q��?             @        ������������������������       �                      @        D       E                     J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        I       J       	            �?      �?             @        ������������������������       �                     �?        K       L                    �?�q�q�?             @        ������������������������       �                     �?        M       N       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     E@        R       S                   �c@�q�q�?             @       ������������������������       �                     @        T       U                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        W       Z                   �]@X�<ݚ�?             "@        X       Y                     P@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        [       ^                   �N@z�G�z�?             @       \       ]                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        `       �       	          ����?�ʍf��?�            �s@       a       �                    �?��<�`�?�            `p@       b       �                   Hp@x!'ǯ�?�            �k@       c       p       
             �?�h:�)�?a            �c@        d       i                    �?
j*D>�?             :@        e       f                    b@r�q��?	             (@        ������������������������       �                     @        g       h       	          ����?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        j       k                   �_@X�Cc�?
             ,@        ������������������������       �                      @        l       o       	          ����?r�q��?             @        m       n                    �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        q       ~       	          pff�?�-�[�?N            ``@       r       }                    �?0x�!���?I            �]@        s       v                    �D@\-��p�?             =@        t       u                   `j@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        w       x                   �c@$�q-�?             :@       ������������������������       �                     3@        y       |                   0f@����X�?             @       z       {                    �E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        7            �V@               �                   @e@�q�q�?             (@       �       �                   `b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ]@�4��?+            @P@        �       �                   �r@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?��h!��?&            �L@        �       �       	          ����?�q�q�?	             .@       ������������������������       �                     "@        �       �                    �L@r�q��?             @        ������������������������       �                     @        �       �                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �g@؇���X�?             E@       �       �       	            �?ףp=
�?             D@       �       �                    �N@`Jj��?             ?@       �       �                   `q@(;L]n�?             >@        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        ������������������������       �                     �?        �       �                    �M@�<ݚ�?             "@        �       �                   xp@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                     K@�G�z��?             D@        �       �                    �?��s����?             5@        �       �                    �H@�����H�?             "@       �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?      �?             (@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   u@�d�����?             3@       �       �                   P`@@�0�!��?             1@       ������������������������       �                     $@        �       �                    @և���X�?             @       �       �       	          ����?z�G�z�?             @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �a@"pc�
�?            �K@       ������������������������       �                     ;@        �       �                    �?X�Cc�?             <@        ������������������������       �                     @        �       �                    e@\X��t�?             7@       �       �                   �c@X�Cc�?	             ,@       �       �       	          `ff�?      �?              @        ������������������������       �                     �?        �       �                    m@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�����H�?             "@       �       �                   �a@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �              
             �?��-�_�?�            0t@       �       �                    �?h�N��?�            pp@       �       �                   @e@x�����?�            �g@        �       �                   �a@P����?%            �M@       ������������������������       �        !             K@        �       �                   `X@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �e@�禺f��?\            �`@        ������������������������       �                     @        �       �       	          ����?     |�?[             `@        �       �                    �?O�o9%�?-            �Q@       �       �                    `@�? Da�?'            �O@        �       �                    @L@�q�q�?             8@       �       �                   �c@�8��8��?
             (@       ������������������������       �        	             &@        ������������������������       �                     �?        �       �                   �X@      �?             (@        ������������������������       �                     @        �       �       	          tff�?      �?              @        ������������������������       �                     @        �       �                   `^@      �?             @        ������������������������       �                     �?        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����? ���J��?            �C@        �       �                   �\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @@        �       �                   0o@      �?              @       �       �                    �H@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �F@���U�?.            �L@        �       �       	             @z�G�z�?             @        ������������������������       �                      @        �       �                    �E@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    @M@ pƵHP�?)             J@       ������������������������       �                     >@        �       �                   q@���7�?             6@       ������������������������       �                     0@        �       �                   `q@r�q��?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    p@�k~X��?+             R@       ������������������������       �                     J@        �       �       	             @P���Q�?             4@       ������������������������       �                     2@        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �G@�0u��A�?#             N@                                hq@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @                                 �?�z�G��?             I@                               �e@� ��1�?            �D@                                �?8�Z$���?            �C@                               �^@���7�?             6@        	      
                  �]@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@                    	          ����?�t����?	             1@                               �r@�q�q�?             (@                               �]@      �?             $@        ������������������������       �                     @                                `_@����X�?             @        ������������������������       �                      @                                �a@���Q��?             @                   	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                 �M@�<ݚ�?             "@       ������������������������       �                     @                                  P@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�b��<     h�h)h,K ��h.��R�(KMKK��hb�B�  S��6�?ם,�d�?�=��!�?b	G��y�?*�Y7�"�?�S�n�?��o��o�?�A�A�?|�W|�W�?�A�A�?      �?        �������?�������?              �?(������?^Cy�5�?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?              �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�?�������?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?      �?                      �?��-��-�?�A�A�?      �?      �?      �?                      �?$��Co�?x�!���?333333�?�������?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?              �?        _^,N��?v����(�?��Q`��?�<�]?[�?Ȥx�L��?�֡�l�?;�;��?;�;��?      �?      �?      �?                      �?      �?      �?'�l��&�?�l��&��?�������?�������?UUUUUU�?UUUUUU�?      �?        y�5���?Cy�5��?�������?�������?۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?        �q�q�?r�q��?      �?      �?              �?      �?        �������?�������?      �?      �?              �?      �?                      �?���?��;���?���*N�?h�T��?7�"�u��?#�u�)��?�,��O�?��O[h��?;�;��?b'vb'v�?UUUUUU�?�������?              �?�������?333333�?              �?      �?        %I�$I��?�m۶m��?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?�[���?qBJ�eD�?��~���?�5�5�?a����?�{a���?UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?;�;��?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?              �?        �R+�R+�?�Z��Z��?      �?      �?              �?      �?        Hp�}�?p�}��?UUUUUU�?UUUUUU�?              �?�������?UUUUUU�?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?�������?�������?���{��?�B!��?�������?�?۶m۶m�?�$I�$I�?              �?      �?              �?                      �?9��8���?�q�q�?      �?      �?              �?      �?              �?                      �?�������?�������?z��y���?�a�a�?�q�q�?�q�q�?      �?      �?              �?      �?              �?              �?      �?      �?      �?      �?                      �?      �?        y�5���?Cy�5��?�������?ZZZZZZ�?              �?۶m۶m�?�$I�$I�?�������?�������?      �?      �?              �?      �?                      �?      �?              �?        F]t�E�?/�袋.�?              �?�m۶m��?%I�$I��?              �?��Moz��?!Y�B�?%I�$I��?�m۶m��?      �?      �?      �?        �$I�$I�?�m۶m��?              �?      �?              �?        �q�q�?�q�q�?�������?�������?              �?      �?                      �?Gb,��o�?n�����?����p�? i��q�?�d�hκ??o��2��?'u_[�?�V'u�?              �?�������?�������?      �?                      �?m��&�l�?e�M6�d�?      �?              �?     @�?��RO�o�?�D+l$�?AA�?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�A�A�?��-��-�?�$I�$I�?۶m۶m�?      �?                      �?              �?      �?      �?�������?UUUUUU�?              �?      �?                      �?p�}��?	�#����?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ;�;��?'vb'vb�?              �?F]t�E�?�.�袋�?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?�q�q�?�8��8��?              �?�������?ffffff�?              �?      �?      �?      �?                      �?�������?�������?�������?�������?      �?                      �?333333�?ffffff�?������?������?;�;��?;�;��?F]t�E�?�.�袋�?      �?      �?              �?      �?                      �?�������?�������?�������?�������?      �?      �?      �?        �$I�$I�?�m۶m��?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?      �?        9��8���?�q�q�?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJv~�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK߅�h��B�7         �       
             �?SH7�j�??           ��@              I                    �?~x�V��?L           �@               H                   f@�+����?�            �k@                                 ``@~��R���?�            �j@                      
             �?$�q-�?(            @P@                                  @^@�z�G��?             $@              
                    �?      �?             @              	                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                   �?h㱪��?"            �K@                                   �Q@8�Z$���?
             *@       ������������������������       �        	             &@        ������������������������       �                      @        ������������������������       �                     E@               '                    �?�����?\            `b@                                  �]@ףp=
�?(             N@        ������������������������       �                     3@                                   �?�p ��?            �D@                                  �a@      �?              @        ������������������������       �                     @                                  pc@z�G�z�?             @        ������������������������       �                     @                      	          033@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                  ``@�FVQ&�?            �@@        ������������������������       �        	             0@                                   @h@�t����?             1@        ������������������������       �                     �?        !       "                    �?      �?             0@        ������������������������       �                     @        #       $       	             �?$�q-�?	             *@       ������������������������       �                     $@        %       &                   �]@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        (       +                    @F@������?4            �U@        )       *                    �B@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ,       5                    �?�s��:��?-             S@        -       4       	          ����?r�q��?             8@       .       3                   pe@      �?	             0@       /       0       	          ����?z�G�z�?             .@        ������������������������       �                     @        1       2                    a@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        6       G       	          ���@R�}e�.�?             J@       7       :       
             �?���c�H�?            �H@        8       9                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ;       F                   ``@�T|n�q�?            �E@       <       E                   Pp@ �o_��?             9@       =       @                    @L@��S���?	             .@        >       ?                     I@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        A       B                    `@      �?              @       ������������������������       �                     @        C       D       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     2@        ������������������������       �                     @        ������������������������       �                     $@        J       Q                   �Z@��&�|�?�            �s@        K       L                   Pa@X�Cc�?	             ,@       ������������������������       �                     @        M       N                   �b@����X�?             @        ������������������������       �                     @        O       P                    �F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        R       }                   `f@���n4s�?�            s@       S       j       	          ����?ཕvt�?�            �r@        T       U                   �i@��Wv��??             [@       ������������������������       �        "            �N@        V       e                   `a@��0{9�?            �G@       W       X                   0j@�+e�X�?             9@        ������������������������       �                      @        Y       \                    �G@�㙢�c�?             7@        Z       [                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ]       ^                   �Y@�����H�?             2@        ������������������������       �                     "@        _       d                    �?�<ݚ�?             "@       `       c       	          433�?      �?              @        a       b       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        f       g                   pb@���7�?             6@        ������������������������       �                     $@        h       i                    �H@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        k       n                    �D@8�o+�?v            �g@        l       m                    i@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        o       t                   8p@�]0��<�?q            �f@       p       s                   �[@ �O�H�?E            �[@        q       r       	          `ff�?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �        @            �X@        u       x                   Xp@�n���?,             R@        v       w                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        y       z                     M@�nkK�?*            @Q@       ������������������������       �                    �F@        {       |                   @b@      �?             8@       ������������������������       �                     5@        ������������������������       �                     @        ~                           �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   @E@T�/�J|�?�            �w@        �       �                    Z@����>�?            �B@        ������������������������       �                      @        �       �                   �]@4�2%ޑ�?            �A@        �       �                   @\@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �       	          hff�?8�Z$���?             :@        �       �                    �?և���X�?             @       �       �                    �?���Q��?             @       �       �                    �L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�}�+r��?             3@       �       �                   c@ףp=
�?	             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    @L@hS>)��?�            @u@       �       �       	          pff�? ��&�?�            �p@       �       �                   �g@������?�             l@       �       �                    �?`��r��?�            �k@        �       �                    �?*
;&���?             G@        ������������������������       �                     &@        �       �                    `@z�G�z�?            �A@       �       �                    �B@�����?             3@        ������������������������       �                      @        �       �                   0c@������?             1@       ������������������������       �                     "@        �       �                     I@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    e@      �?
             0@       ������������������������       �        	             .@        ������������������������       �                     �?        �       �                   @[@�O"9��?t             f@        �       �                   `m@      �?              @       ������������������������       �                     @        �       �                   `d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        m             e@        ������������������������       �                     �?        �       �                    `@d}h���?             E@        �       �                   �f@      �?             (@        ������������������������       �                     @        �       �                    @I@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                    @K@ףp=
�?             >@       �       �                    o@ 	��p�?             =@       ������������������������       �                     8@        �       �                   `a@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `f@���+�?0            �R@        �       �                   @_@�q�q�?             "@        ������������������������       �                     @        �       �                   �b@      �?             @        ������������������������       �                      @        �       �                   �d@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    ]@�θ�?+            @P@        �       �                    �?����X�?             @       ������������������������       �                     @        �       �                   0p@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @M@д>��C�?&             M@        �       �                   �t@X�<ݚ�?             "@       �       �                   0n@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �r@ i���t�?            �H@       �       �                    b@P�Lt�<�?             C@       ������������������������       �                     :@        �       �                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   �c@���|���?             &@       �       �                   �`@�q�q�?             @        ������������������������       �                      @        �       �                     O@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   @t@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ���t��?�~�E)�?���X�?VR�{���?�+c���?jNq��?�[�琚�?R����?;�;��?�؉�؉�?333333�?ffffff�?      �?      �?      �?      �?              �?      �?                      �?              �?��)A��?־a���?;�;��?;�;��?              �?      �?                      �?q�{���?G-B���?�������?�������?              �?��+Q��?Q��+Q�?      �?      �?      �?        �������?�������?              �?      �?      �?      �?                      �?|���?>����?              �?�?<<<<<<�?      �?              �?      �?              �?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?              �?      �?        J��/�?m��֡�?]t�E�?F]t�E�?              �?      �?        �k(���?��k(��?�������?UUUUUU�?      �?      �?�������?�������?      �?              �?      �?      �?                      �?              �?      �?        �;�;�?'vb'vb�?/�����?4և����?UUUUUU�?UUUUUU�?      �?                      �?6eMYS��?���)k��?�Q����?
ףp=
�?�������?�?۶m۶m�?�$I�$I�?              �?      �?              �?      �?              �?      �?      �?              �?      �?                      �?              �?      �?              �?        ��9Hڰ?������?�m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ^���۪?��xAR�?����?.�$�?{	�%���?�^B{	��?              �?L� &W�?m�w6�;�?���Q��?R���Q�?      �?        d!Y�B�?�7��Mo�?�������?333333�?      �?                      �?�q�q�?�q�q�?              �?�q�q�?9��8���?      �?      �?      �?      �?              �?      �?                      �?      �?        F]t�E�?�.�袋�?              �?UUUUUU�?UUUUUU�?      �?                      �?�-q��ܢ?#�X�0��?�$I�$I�?۶m۶m�?      �?                      �?;ڼOqɠ?\2�h��?5'��Ps�?c��2��?UUUUUU�?UUUUUU�?      �?                      �?              �?r�qǱ?r�q��?UUUUUU�?UUUUUU�?              �?      �?        d!Y�B�?�Mozӛ�?              �?      �?      �?              �?      �?        �$I�$I�?�m۶m��?              �?      �?        gq�T�e�?f:z��h�?���L�?�u�)�Y�?      �?        �A�A�?�������?�q�q�?r�q��?              �?      �?        ;�;��?;�;��?۶m۶m�?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?(�����?�5��P�?�������?�������?              �?      �?                      �?TTTTTT�?]]]]]]�?Z�iu���?,�T�R�?n۶m۶�?%I�$I��?������?�p"^�?���,d!�?8��Moz�?      �?        �������?�������?Q^Cy��?^Cy�5�?              �?xxxxxx�?�?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?Cr����?��F($w?      �?      �?      �?              �?      �?              �?      �?              �?                      �?I�$I�$�?۶m۶m�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?������?�{a���?      �?        333333�?�������?      �?                      �?              �?�n0E>��?�"�u�)�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?              �?      �?        ى�؉��?�؉�؉�?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?a���{�?|a���?�q�q�?r�q��?UUUUUU�?�������?      �?                      �?      �?        /�����?����X�?���k(�?(�����?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJwm�ohG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@>         �       
             �?<qn�h��?=           ��@              O                    �?0��k���?F           @�@              
                   �Z@_n8�?�            �u@               	                    �?�q�q�?             (@                                   �?r�q��?             @        ������������������������       �                     @                      	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @               $                    �?t�e�í�?�            �t@                                  �`@p�ݯ��?             C@                                   �O@ҳ�wY;�?             1@                     
             �?և���X�?             ,@        ������������������������       �                     �?                                  @[@�n_Y�K�?
             *@        ������������������������       �                      @                                    F@���!pc�?             &@        ������������������������       �                     �?                                   �?z�G�z�?             $@                                  �?�����H�?             "@        ������������������������       �                     @                                   `@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               #                    b@؇���X�?             5@                       	          ����?և���X�?             @                                   �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        !       "       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        %       8                    �? 7���B�?�            �r@       &       /       	          ����? '�Ӕ�?�            �j@        '       (                   �g@��<D�m�?#            �H@        ������������������������       �                     5@        )       *       	          ����? �Cc}�?             <@       ������������������������       �                     8@        +       .                   �_@      �?             @        ,       -                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        0       1                   �Q@�dJ�Ҙ?k            `d@        ������������������������       �                     �?        2       3                   @s@ A��� �?j            @d@       ������������������������       �        Z            �a@        4       7       
             �?���N8�?             5@        5       6                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     2@        9       N       	          ����?p��@���?0            @U@       :       ;                   �[@��2(&�?             F@        ������������������������       �                     �?        <       A                   �i@X�EQ]N�?            �E@       =       @                   �_@XB���?             =@        >       ?                   �^@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     6@        B       K                   �_@����X�?	             ,@       C       D                   �_@ףp=
�?             $@        ������������������������       �                     @        E       J                    �?r�q��?             @       F       I                   �a@      �?             @        G       H                     P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        L       M       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �D@        P       }                   �b@F�H~4o�?f            �e@       Q       \                    �?����X��?D             \@        R       S       
             �?��Q��?
             4@        ������������������������       �                     �?        T       [       	          ����?p�ݯ��?	             3@       U       X                    @L@�q�q�?             (@       V       W                    ]@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        Y       Z                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ]       ^                   @Y@�3Ea�$�?:             W@        ������������������������       �                      @        _       b                    @F@:	��ʵ�?9            �V@        `       a                    W@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        c       t                   pb@�����	�?6            @U@       d       o       	          033�?��a�n`�?(             O@        e       j                    @K@�GN�z�?             6@        f       i                   Pa@X�<ݚ�?             "@       g       h                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        k       n                    �?$�q-�?	             *@        l       m                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        p       q                   �b@�(\����?             D@       ������������������������       �                    �B@        r       s       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        u       v                   �_@��+7��?             7@        ������������������������       �                     &@        w       z                    �?      �?             (@       x       y                   @b@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        {       |                    �L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                    �H@�'N��?"            �N@               �                    �F@�f7�z�?             =@       �       �                    �?@�0�!��?	             1@       �       �       	          ����?@4և���?             ,@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �       �       	          033@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             (@        �       �       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?     ��?             @@        ������������������������       �                     (@        �       �       
             �?      �?             4@        ������������������������       �                     @        �       �                    p@�q�q�?	             .@       �       �                   @W@r�q��?             (@        �       �                    �N@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�y���?�            �x@       �       �                    �?��� �6�?�            �t@       �       �                    �?�S=ث?�?�            r@        �       �                    q@ڡR����?            �H@       �       �       	          ����?      �?             <@       �       �       	             �?�C��2(�?             6@       �       �                   pd@�����?             5@        ������������������������       �                     @        �       �                   @n@؇���X�?	             ,@       �       �                   @k@�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   Pe@�ՙ/�?
             5@       �       �                    �K@�q�q�?             (@       �       �       	          @33�?      �?              @        �       �                   0d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @G@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?�             n@        �       �                    b@�2����?!            �K@       �       �                   �Y@ףp=
�?             I@        �       �                   �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �I@���.�6�?             G@       ������������������������       �                     <@        �       �                    @J@r�q��?
             2@        ������������������������       �                      @        �       �                    X@      �?	             0@        �       �       	          @33�?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        �       �                   �b@z�G�z�?             @        ������������������������       �                      @        �       �                   `m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?f�1�?p             g@       ������������������������       �        :            �X@        �       �                   �c@ 	��p�?6            �U@       �       �                   �b@H%u��?             I@       �       �                    �?`Ӹ����?            �F@        �       �                   �^@�t����?             1@        �       �                    ^@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     <@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �B@        �       �                    V@և���X�?             E@        ������������������������       �        
             1@        �       �                   @`@`2U0*��?             9@        �       �       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �       �                    �?�2�,��?*            �P@       �       �                    �?��C���?            �G@       �       �                    �?d��0u��?             >@        ������������������������       �                     @        �       �                   �]@l��
I��?             ;@        �       �                    Z@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   pf@R���Q�?             4@       �       �                   `W@�KM�]�?             3@        �       �                   �_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �        
             1@        �       �                    �G@�z�G��?             4@        ������������������������       �                     @        �       �                   @n@      �?
             0@       ������������������������       �                      @        �       �                   �`@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �g�g�?!�v!�v�?��؉���?�؉�؉�?�����!�?B�`�;�?�������?�������?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�rv��?�1����?Cy�5��?^Cy�5�?�������?�������?�$I�$I�?۶m۶m�?              �?;�;��?ى�؉��?              �?F]t�E�?t�E]t�?              �?�������?�������?�q�q�?�q�q�?      �?              �?      �?              �?      �?                      �?      �?        �$I�$I�?۶m۶m�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?h/�����?	�%����?�V�9�&�?HM0��>�?և���X�?��S�r
�?              �?۶m۶m�?%I�$I��?              �?      �?      �?      �?      �?      �?                      �?      �?        )��I� �?w��|��?      �?        �����Hy?,R�n��?              �?�a�a�?��y��y�?UUUUUU�?UUUUUU�?              �?      �?                      �?�?�������?t�E]t�?��.���?      �?        qG�wĽ?w�qG�?�{a���?GX�i���?�$I�$I�?۶m۶m�?              �?      �?                      �?�$I�$I�?�m۶m��?�������?�������?              �?UUUUUU�?�������?      �?      �?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?                      �?u�g���?F5�� �?n۶m۶�?I�$I�$�?�������?ffffff�?      �?        ^Cy�5�?Cy�5��?�������?�������?�$I�$I�?۶m۶m�?      �?                      �?�������?�������?      �?                      �?      �?        ��,d!�?����7��?      �?        l�l��?��O��O�?�������?�������?              �?      �?        �?{{{{{{�?�c�1Ƹ?�s�9��?]t�E�?�袋.��?�q�q�?r�q��?�$I�$I�?�m۶m��?              �?      �?              �?        ;�;��?�؉�؉�?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?Y�B��?zӛ����?              �?      �?      �?�$I�$I�?�m۶m��?      �?                      �?�������?�������?              �?      �?        �����?ާ�d��?O#,�4��?a���{�?ZZZZZZ�?�������?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?�큍��?
H�Ʌ��?)�k?J��?\�Q�~�?�.k���?j���� �?����S��?����X�?      �?      �?]t�E�?F]t�E�?=��<���?�a�a�?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?      �?              �?        UUUUUU�?�������?              �?      �?        �a�a�?�<��<��?�������?�������?      �?      �?      �?      �?              �?      �?              �?                      �?�q�q�?�q�q�?      �?                      �?      �?      �?��7�}��?� O	��?�������?�������?      �?      �?      �?                      �?���7���?Y�B��?      �?        �������?UUUUUU�?              �?      �?      �?      �?      �?      �?                      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        e�kBP��?�	A����?      �?        ������?�{a���?)\���(�?���Q��??�>��?l�l��?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?�������?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?���Q��?{�G�z�?      �?      �?      �?                      �?      �?        o�Wc"=�?"=P9���?L� &W�?g���Q��?wwwwww�?DDDDDD�?      �?        h/�����?Lh/����?�m۶m��?�$I�$I�?              �?      �?        333333�?333333�?(�����?�k(���?      �?      �?      �?                      �?              �?      �?              �?        333333�?ffffff�?      �?              �?      �?              �?      �?      �?              �?      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$ֽQhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@A         p       	          ����?TU�`��?<           ��@              E                    �?(b>+��?$           P}@                      
             �?��"���?z            @i@               	                   �k@<����?=            �W@                     	          ����? _�@�Y�?&             M@       ������������������������       �        !            �J@                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        
                           �?��G���?            �B@                                  �?�q�q�?             8@                                  �?�GN�z�?             6@                                   �?�z�G��?             $@        ������������������������       �                      @                                  @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                   _@r�q��?             (@        ������������������������       �                     @                                  0a@�q�q�?             @                                  �I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@               "                    P@xZ�l ��?=            �Z@               !                    �?�t����?             1@                                   �?r�q��?             (@                      	          @33�?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        #       >                    @M@>���a��?2            �V@       $       /                   `\@      �?+             T@        %       *                    �?�q�q�?             2@        &       '                   �_@և���X�?             @        ������������������������       �                      @        (       )                    �G@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        +       ,                   �b@"pc�
�?             &@       ������������������������       �                     @        -       .                   �k@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        0       1                   �k@`Jj��?             O@        ������������������������       �        	             3@        2       5                    l@�ʈD��?            �E@        3       4                    a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        6       =                   ``@�7��?            �C@        7       <                   �r@�����?
             5@       8       ;                   �q@r�q��?             (@       9       :                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        
             2@        ?       D                    �?�z�G��?             $@       @       C                    b@      �?             @       A       B                   Hq@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        F       I                   �O@V#L��?�            �p@        G       H       
             �?`�Q��?             9@       ������������������������       �        
             1@        ������������������������       �                      @        J       k                    c@�R����?�            @n@       K       N                   �W@$�q-�?�            �k@        L       M                   �V@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        O       b       
             �?��}$�6�?�            �j@        P       [       	          ����?���Q��?             >@       Q       Z                    g@����X�?             ,@       R       Y                    �?�θ�?             *@        S       T                    �?      �?             @        ������������������������       �                      @        U       X                   �`@      �?             @        V       W                   `l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        \       a                    �?      �?             0@       ]       `                   �b@��S�ۿ?             .@        ^       _                    �K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        c       j                    �?��W��#�?x             g@        d       i                    �?��v$���?*            �N@        e       f                   �r@�8��8��?	             (@       ������������������������       �                     $@        g       h                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        !            �H@        ������������������������       �        N            �^@        l       m                    �K@�q�q�?             5@       ������������������������       �                     (@        n       o                    �N@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        q       �                   �b@*�h�.Z�?           |@       r       �                    �?j\4F��?�            �w@        s       �                    �?�ĚpF�?4            @U@       t       �                    �?*;L]n�?#             N@       u       �                    �?�n_Y�K�?             J@        v       y                   @p@�E��ӭ�?
             2@        w       x                   �\@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        z       {       	          ����?      �?              @        ������������������������       �                     @        |       }       	             �?z�G�z�?             @        ������������������������       �                     �?        ~                          �a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?H�V�e��?             A@        ������������������������       �                     @        �       �                    `@��� ��?             ?@        ������������������������       �                     .@        �       �       	          ����?      �?             0@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `c@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                    a@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?HP�s��?             9@        �       �                   @Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Xw@���7�?             6@       ������������������������       �                     5@        ������������������������       �                     �?        �       �                   �[@ؓFl:8�?�            Pr@        �       �                    �?     ��?             @@       �       �                   `_@�<ݚ�?             ;@        ������������������������       �                     .@        �       �                    �?      �?             (@       �       �       	          033@���Q��?             $@       �       �                   0b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   P`@4��6�?�            Pp@        �       �                    �?\�ih�<�?6            �W@        ������������������������       �                     6@        �       �       	          ����?z�z�7��?*            @R@        �       �                    �G@��X��?             <@        ������������������������       �                     @        �       �                    �?�û��|�?             7@       �       �                   0p@      �?	             0@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@       �       �                   @s@�����H�?             "@        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �q@؇���X�?             @        ������������������������       �                     @        �       �                    [@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �I@�:�^���?            �F@        ������������������������       �                     .@        �       �                   h@�r����?             >@        �       �       	             �?���Q��?             $@        �       �                    �?���Q��?             @       �       �                    @K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `^@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        �       �       
             �?x�}���?i            �d@        �       �                   �c@�<ݚ�?             2@       ������������������������       �                     $@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   �e@PL��V�?]            �b@       �       �       	          ����?��[����?U             a@        �       �                    �?��?^�k�?            �A@        ������������������������       �                     2@        �       �                   @b@�IєX�?             1@       ������������������������       �                     &@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        B            �Y@        �       �                     L@"pc�
�?             &@        ������������������������       �                     @        �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   Xr@`��_��?4            �Q@       �       �                   �o@l`N���?(            �J@       �       �                    �?�p ��?!            �D@        �       �                    �?z�G�z�?             .@        �       �       	          033�?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �F@�C��2(�?	             &@        �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �       	             @�	j*D�?             :@       �       �       
             �?@�0�!��?             1@        ������������������������       �                     �?        �       �                   �i@      �?             0@        �       �                    e@      �?             @       �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             (@        �       �                    `@X�<ݚ�?             "@        ������������������������       �                     @        �       �                    W@�q�q�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �             	          ���@�<ݚ�?             2@       �       �                   c@@�0�!��?             1@        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �I@@4և���?	             ,@                                �r@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��hb�BP  ��Fc*�?y�\���?�N�I�?%�b�l��?�2|#
L�?��A����?�X�0Ҏ�?���%N�?�{a���?#,�4�r�?              �?�������?�������?      �?                      �?v�)�Y7�?#�u�)��?�������?�������?]t�E�?�袋.��?333333�?ffffff�?      �?              �?      �?      �?                      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�w�Zn�?�+J�#�?�?<<<<<<�?UUUUUU�?�������?�������?333333�?      �?                      �?              �?              �?J��I���?؂-؂-�?      �?      �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?        /�袋.�?F]t�E�?      �?        333333�?�������?      �?                      �?���{��?�B!��?      �?        A_���?�}A_з?      �?      �?      �?                      �?��[��[�?�A�A�?=��<���?�a�a�?�������?UUUUUU�?]t�E�?F]t�E�?      �?                      �?              �?      �?              �?        333333�?ffffff�?      �?      �?      �?      �?      �?                      �?              �?              �?�5Xl�?:)�Nʧ�?{�G�z�?��(\���?              �?      �?        �������?���!pc�?�؉�؉�?;�;��?۶m۶m�?�$I�$I�?      �?                      �?M�w�Z�?7��XQ�?333333�?�������?�$I�$I�?�m۶m��?�؉�؉�?ى�؉��?      �?      �?              �?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?              �?      �?�������?�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?��Moz��?d!Y�Bv?.�u�y�?;ڼOqɐ?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?      �?        �q�q�?9��8���?              �?      �?        �F��?>S�޹:�?�?�����?�V�Z�?�?uuuuuu�?�������?""""""�?ى�؉��?;�;��?�q�q�?r�q��?�������?�������?              �?      �?              �?      �?              �?�������?�������?      �?              �?      �?      �?                      �?ZZZZZZ�?iiiiii�?      �?        �B!��?�{����?              �?      �?      �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?{�G�z�?q=
ףp�?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?�.�袋�?              �?      �?        Y���?ܴE��?      �?      �?�q�q�?9��8���?              �?      �?      �?333333�?�������?�������?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?      �?        Q��kꝳ?�n��B��?Ai�
��?�%N���?              �?�lٲe��?ҤI�&M�?%I�$I��?n۶m۶�?              �?��,d!�?8��Moz�?      �?      �?              �?�������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?        l�l��?}�'}�'�?              �?�?�������?�������?333333�?333333�?�������?      �?      �?      �?                      �?              �?�������?�������?              �?      �?                      �?4u~�!��?�(፦�?�q�q�?9��8���?              �?      �?      �?              �?      �?        L�Ϻ��?�u�)�Y�?������}?�8R4��?�A�A�?_�_��?              �?�?�?              �?UUUUUU�?�������?              �?      �?                      �?F]t�E�?/�袋.�?              �?�$I�$I�?�m۶m��?              �?      �?        6��9�?��ۥ���?
�[���?�R���?dp>�c�?8��18�?�������?�������?      �?      �?              �?      �?        F]t�E�?]t�E�?      �?      �?      �?                      �?              �?vb'vb'�?;�;��?ZZZZZZ�?�������?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �q�q�?r�q��?              �?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        9��8���?�q�q�?ZZZZZZ�?�������?UUUUUU�?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?�������?�������?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�[KhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�@         �                    �?�m=62}�?B           ��@              +                    `@�p�*��?[           Ё@                                   �?�!�z�0�?<            �Z@                                  �?      �?&             P@                                   �O@�㙢�c�?             7@                                 �Z@��2(&�?             6@        ������������������������       �                     �?                                   �?�����?             5@       	       
                    �?�r����?
             .@        ������������������������       �                      @                                    J@8�Z$���?	             *@        ������������������������       �                     �?                                  �`@�8��8��?             (@       ������������������������       �                     "@                                  pb@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �D@               &       	          hff @�&!��?            �E@                     
             �?�g�y��?             ?@                                  `Q@�q�q�?	             2@                     
             �?؇���X�?             ,@        ������������������������       �                     �?                                   @$�q-�?             *@                                 �X@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @                %                   `@�θ�?             *@        !       "                    �?      �?             @        ������������������������       �                      @        #       $       	             п      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        '       (                    �?�8��8��?             (@        ������������������������       �                      @        )       *       	          `ff@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ,       q       
             �?�b��z�?           �|@        -       `                   �o@��!L:A�?c            �d@       .       ?                    �?X��ʑ��?:            �U@        /       >       	          `ff@��a�n`�?             ?@       0       3                    �?д>��C�?             =@        1       2                   �a@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        4       ;                   0e@������?             1@       5       6       	          ����?؇���X�?	             ,@        ������������������������       �                     @        7       :                    �H@      �?              @        8       9                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        <       =                   `^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        @       K                    �?��N`.�?(            �K@        A       J                    �N@     ��?
             0@       B       I                   �`@�eP*L��?             &@       C       D                   �\@      �?              @        ������������������������       �                     �?        E       F                   �_@؇���X�?             @        ������������������������       �                     @        G       H                    �K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        L       _                    �?:�&���?            �C@       M       X                   �a@��a�n`�?             ?@       N       S                    j@ףp=
�?             4@        O       R                    �E@z�G�z�?             @       P       Q                   pg@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       U                    �O@��S�ۿ?
             .@       ������������������������       �                     *@        V       W                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z       	          ����?�eP*L��?
             &@        ������������������������       �                     @        [       \                     G@����X�?             @        ������������������������       �                     @        ]       ^                   Pc@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        a       h                   �r@���R�?)            @T@       b       c                    �I@�X�C�?             L@        ������������������������       �        
             1@        d       e                   pa@�θ�?            �C@        ������������������������       �                     4@        f       g                    �M@�\��N��?
             3@        ������������������������       �                     "@        ������������������������       �                     $@        i       j                   �s@�q�����?             9@        ������������������������       �                     "@        k       p       	          ����?      �?
             0@       l       o                     L@և���X�?             @        m       n                    e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        r       u                    c@�L���?�            �r@        s       t                   �b@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        v       �                   �g@��� @�?�            r@       w       �                   �r@�n���?�             r@       x       y                    �?8�M'��?�            �m@        ������������������������       �        1            �R@        z       �                    @L@c��3�?i            @d@       {       �                   �[@ ���z��?R            �_@        |       �                   �c@      �?             0@       }       �                    �?�<ݚ�?             "@       ~       �                    �?      �?              @               �                     D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        F            �[@        �       �                    @��R[s�?            �A@       �       �                    �L@r�q��?             >@        �       �                   �a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?HP�s��?             9@        ������������������������       �                     "@        �       �       	             �?      �?             0@       �       �                    b@��S�ۿ?
             .@       ������������������������       �                     *@        �       �                   P`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    a@z�G�z�?             @        ������������������������       �                     @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �L@@�0�!��?            �I@       ������������������������       �                     >@        �       �                   pe@և���X�?
             5@       �       �                    �?��.k���?	             1@       �       �       	          @33�?�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �u@����X�?             @        �       �                     O@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �b@�=C|F�?�            �u@       �       �                   Pf@ܾ�z�<�?�            �s@        �       �                   @^@�]���?I            �\@        �       �       
             �?P���Q�?             D@       ������������������������       �                     >@        �       �                   �\@z�G�z�?             $@        ������������������������       �                     @        �       �                    a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        0            �R@        �       �       	          ����?0sS]�?�            �h@        �       �                    �?&�a2o��?3            @Q@        �       �       	          hff�?�8��8��?             8@       �       �       
             �?r�q��?	             (@       ������������������������       �                     "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        �       �       
             �?f.i��n�?"            �F@       �       �       	          ����?x�����?            �C@        ������������������������       �                     *@        �       �                    @L@�	j*D�?             :@       �       �                    �?      �?             0@       �       �                    b@��S�ۿ?
             .@       ������������������������       �                     "@        �       �                    �?r�q��?             @       �       �                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �q@���Q��?             $@        �       �                   �[@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    w@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �R@     ��?R             `@       �       �                    �J@�&/�E�?P             _@        �       �                    �?8�Z$���?            �C@       �       �                    �I@�#-���?            �A@       ������������������������       �                     8@        �       �                   �`@���!pc�?             &@       �       �                    @J@�����H�?             "@       ������������������������       �                     @        �       �                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	             @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ����?`��>�ϗ?9            @U@        �       �                     P@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �        2            @R@        �       �       	             @      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @G@)O���?             B@        �       �                   �f@      �?             (@       �       �                    `@ףp=
�?             $@       �       �                    @D@r�q��?             @        �       �                    �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   c@�q�q�?             8@        ������������������������       �                      @        �                          �M@���!pc�?             6@       �       �                    a@և���X�?             ,@        �       �                    d@r�q��?             @        ������������������������       �                     @        �       �       	          @33�?�q�q�?             @       �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     M@      �?              @       ������������������������       �                     @                                 �h@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �t�b�]     h�h)h,K ��h.��R�(KMKK��hb�B0  ��f���?w>�̓�?�@i�
�?�~�-q��?��XQ�?�ީk9��?      �?      �?d!Y�B�?�7��Mo�?t�E]t�?��.���?      �?        �a�a�?=��<���?�?�������?              �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?S֔5eM�?֔5eMY�?�B!��?��{���?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?�������?�������?      �?                      �?              �?      �?        ى�؉��?�؉�؉�?      �?      �?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        J�nH�8�?m�"o��?J�����?�'����?��}A�?�}A_�?�c�1��?�s�9��?a���{�?|a���?UUUUUU�?UUUUUU�?      �?                      �?xxxxxx�?�?۶m۶m�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?� O	��?��oX���?      �?      �?t�E]t�?]t�E�?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �o��o��?�A�A�?�s�9��?�c�1��?�������?�������?�������?�������?      �?      �?              �?      �?                      �?�?�������?              �?      �?      �?              �?      �?        ]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?              �?��ӭ�a�?�)O�?%I�$I��?�m۶m��?              �?�؉�؉�?ى�؉��?              �?�5��P�?y�5���?      �?                      �?�p=
ף�?���Q��?      �?              �?      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?                      �?}���g�?L�Ϻ��?�$I�$I�?۶m۶m�?      �?                      �?���ʻ��?@�0�!��?r�q��?r�qǱ?]��ǃ�?2�N��ç?      �?        �E����?��ӭ�a�?�����~�?�@ �?      �?      �?9��8���?�q�q�?      �?      �?      �?      �?      �?                      �?      �?                      �?      �?              �?        X|�W|��?PuPu�?�������?UUUUUU�?�������?333333�?      �?                      �?q=
ףp�?{�G�z�?      �?              �?      �?�������?�?      �?              �?      �?      �?                      �?              �?�������?�������?              �?      �?      �?      �?                      �?ZZZZZZ�?�������?      �?        �$I�$I�?۶m۶m�?�?�������?333333�?ffffff�?              �?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?J��/�?�C��:��?vb'vb'�?�;�;�?���ϑ?��ʇq�?�������?ffffff�?              �?�������?�������?              �?�������?333333�?      �?                      �?              �?q�)`>�?����g��?ہ�v`��?��Q�g��?UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�>�>��?�`�`�?�A�A�?��o��o�?              �?;�;��?vb'vb'�?      �?      �?�?�������?              �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        333333�?�������?�������?333333�?      �?                      �?�������?�������?      �?                      �?      �?              �?     ��?�s�9�?2�c�1�?;�;��?;�;��?_�_�?�A�A�?              �?t�E]t�?F]t�E�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?      �?                      �?�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?��8��8�?9��8���?      �?      �?�������?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?        t�E]t�?F]t�E�?۶m۶m�?�$I�$I�?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�-�`hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�G         v                   �`@Ly�'^��?A           ��@               7       	          ����?��\m�~�?�             y@               .                    �?�&���?`             c@                                 �T@x>ԛ/��?K            �^@                                   �?�FVQ&�?            �@@                      	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        	       
                    [@�g�y��?             ?@       ������������������������       �                     0@                      
             �?��S�ۿ?	             .@       ������������������������       �                     *@                                    E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �F@���?5            @V@        ������������������������       �        
             6@                                  0i@�d�K���?+            �P@                                  �^@�t����?
             1@       ������������������������       �                     (@                                   �G@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @               #                    �?      �?!             I@                                  �?�q�q�?             8@                                  �`@և���X�?             @                     	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @                                    �?@�0�!��?             1@        ������������������������       �                     @        !       "       
             �?      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        $       +                   �[@�	j*D�?             :@        %       &                   `k@���|���?             &@        ������������������������       �                     @        '       *       	          ����?      �?              @        (       )                   �Y@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ,       -                   �q@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        /       0                    �G@��a�n`�?             ?@        ������������������������       �                     �?        1       6                    @��S�ۿ?             >@       2       3                   @V@XB���?             =@       ������������������������       �                     4@        4       5                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        8       K                    �?�TG!u�?�            �n@        9       J                    `P@և���X�?             5@       :       E                   �q@�t����?             1@       ;       >                    �?r�q��?             (@        <       =                     M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ?       D                    @N@ףp=
�?             $@       @       A                   @_@      �?             @        ������������������������       �                      @        B       C       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        F       I                   �]@���Q��?             @       G       H       	          033�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        L       s                    �Q@@�s��?�            @l@       M       V       
             �?�V���?�            �j@        N       U                   (w@\-��p�?             =@       O       T                    �?�>����?             ;@        P       S                   @^@�q�q�?             @       Q       R                   �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                      @        W       h                    �?�F�sɪ?r            @g@       X       g       	          ����? ���z��?L            �_@       Y       Z                   `_@�g�y��?(             O@       ������������������������       �                     H@        [       ^                   �\@؇���X�?             ,@        \       ]       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        _       `                    �?�8��8��?	             (@        ������������������������       �                     @        a       b       	          ����?      �?              @        ������������������������       �                     �?        c       f                    �F@؇���X�?             @        d       e                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        $            @P@        i       l                    �J@����˵�?&            �M@        j       k                   �_@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        m       r                    X@@�E�x�?            �H@        n       o                    �?؇���X�?             @        ������������������������       �                     @        p       q                     N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     E@        t       u                   �c@�eP*L��?             &@       ������������������������       �                     @        ������������������������       �                     @        w       �       
             �?X�Cc�?J           0�@        x       �                   `a@�q�q�?�            �i@       y       �                    �?     ��?W             `@       z       {                   �U@�θ�?,            @P@        ������������������������       �                     @        |       }                   �e@�n`���?+             O@        ������������������������       �        	             ,@        ~       �                    �M@      �?"             H@              �                    a@     ��?             @@       �       �                   �`@�z�G��?             >@       �       �                   �a@��X��?             <@        �       �                   �h@X�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     M@���y4F�?             3@       �       �                    @G@      �?             0@        �       �                   �r@����X�?             @       �       �                   �b@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �       	          @33�?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �^@      �?	             0@        �       �                    d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        �       �                   �Q@�q�q�?+            �O@        ������������������������       �                     @        �       �                    �K@�d�����?'            �L@       �       �                    �?�KM�]�?             C@       �       �                    �?�L���?            �B@       �       �                    �?Pa�	�?            �@@        �       �                    @D@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     7@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                     H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   `l@D�n�3�?             3@        �       �       	          ����?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�θ�?	             *@        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �L@ףp=
�?             $@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��r�Z}�?/            �S@       �       �       	          ����?`2U0*��?             I@        �       �                    �J@����X�?             @        ������������������������       �                     @        �       �                   �b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �E@        �       �                   �e@J�8���?             =@       �       �                   �j@�+e�X�?             9@        ������������������������       �                     $@        �       �                    �?���Q��?             .@        ������������������������       �                     @        �       �       
             �?"pc�
�?	             &@        ������������������������       �                     �?        �       �                   �l@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                    �?FC�H�k�?�            ps@        �       �       	          033@@9G��?8            �X@       �       �                    �?@��8��?7             X@        �       �                   Pc@$�q-�?             :@        �       �                   �b@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    e@P���Q�?	             4@       ������������������������       �                     ,@        �       �                   �r@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        )            �Q@        ������������������������       �                      @        �       �                    I@Jd+����?�            �j@        �       �                   �`@"pc�
�?             6@        ������������������������       �                      @        �       �                   0f@ףp=
�?             4@       �       �                    �?�X�<ݺ?             2@       �       �                     P@@4և���?
             ,@       ������������������������       �                     &@        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                          �?�Ę�;�?}            �g@        �       �                   �n@��Hg���?            �F@       �       �                   �a@     ��?             @@        ������������������������       �                     (@        �       �                   �k@R���Q�?             4@       �       �                   g@@4և���?             ,@        ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	             @�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �D@�n_Y�K�?             *@        �       �                   �^@      �?             @        ������������������������       �                      @        �       �                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   Pc@�<ݚ�?             "@        ������������������������       �                     @        �                          �?���Q��?             @       �                          f@      �?             @        ������������������������       �                      @                                 @L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                 �L@����1�?c            @b@                                �G@`�c�г?U             _@       ������������������������       �        +            @P@                                 �?�U�:��?*            �M@       	                         �?�q��/��?#             G@       
                        `l@������?             B@       ������������������������       �                     5@                                 m@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@                    	             �?���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@                                �e@8�A�0��?             6@        ������������������������       �                     @                                �\@�\��N��?             3@        ������������������������       �                     @                                 b@      �?
             0@                   	          033�?"pc�
�?             &@                               @f@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?                                  N@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��hb�B�  ȫ�rV��?���T8�?��Q��?���Q��?\�\��?R��Q���?;ڼOq��?�K�`m�?|���?>����?      �?      �?              �?      �?        �B!��?��{���?              �?�?�������?              �?      �?      �?      �?                      �?e%+Y�J�?7��Mmj�?      �?        �rv��?����?<<<<<<�?�?      �?        333333�?�������?              �?      �?              �?      �?�������?�������?۶m۶m�?�$I�$I�?�������?�������?              �?      �?              �?        ZZZZZZ�?�������?      �?              �?      �?              �?      �?        ;�;��?vb'vb'�?]t�E]�?F]t�E�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �?�������?              �?      �?        �c�1Ƹ?�s�9��?      �?        �?�������?�{a���?GX�i���?              �?�q�q�?�q�q�?      �?                      �?      �?        �����߸?@�O%��?۶m۶m�?�$I�$I�?�������?�������?UUUUUU�?�������?      �?      �?      �?                      �?�������?�������?      �?      �?              �?      �?      �?      �?                      �?              �?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        ��	���?��~H��?��V!�n�?D��=��?�{a���?a����?h/�����?�Kh/��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �n�ᆛ?$�<��#�?�@ �?�����~�?�B!��?��{���?              �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?��/���?W'u_�?�������?�������?      �?                      �?9/���?և���X�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?t�E]t�?]t�E�?              �?      �?        %I�$I��?�m۶m��?UUUUUU�?UUUUUU�?     ��?     ��?�؉�؉�?ى�؉��?      �?        �c�1��?�9�s��?              �?      �?      �?      �?      �?333333�?ffffff�?%I�$I��?n۶m۶�?r�q��?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?(������?6��P^C�?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?Cy�5��?y�5���?�k(���?(�����?}���g�?L�Ϻ��?|���?|���?�������?�������?              �?      �?              �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?(������?l(�����?�������?UUUUUU�?              �?      �?        �؉�؉�?ى�؉��?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?      �?                      �?              �?�&��jq�?G�D�#�?{�G�z�?���Q��?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?|a���?�rO#,��?���Q��?R���Q�?              �?�������?333333�?      �?        F]t�E�?/�袋.�?      �?        �������?�������?      �?                      �?      �?        �Σ�)�?��p�X�?������?9/���?UUUUUU�?UUUUUU�?�؉�؉�?;�;��?�������?UUUUUU�?      �?                      �?ffffff�?�������?      �?        �������?UUUUUU�?      �?                      �?      �?                      �?��PI7��?���"��?F]t�E�?/�袋.�?      �?        �������?�������?�q�q�?��8��8�?�$I�$I�?n۶m۶�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?K8����?��W��?؂-؂-�?��I��I�?      �?      �?      �?        333333�?333333�?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?ى�؉��?;�;��?      �?      �?      �?              �?      �?              �?      �?        �q�q�?9��8���?              �?�������?333333�?      �?      �?              �?      �?      �?              �?      �?              �?        �Ν;w��?Ĉ#F��?��Zk���?��RJ)��?      �?        �A�I�?�pR�屵?�B����?��Mozӻ?�q�q�?�q�q�?      �?        �������?�?              �?      �?        333333�?�������?      �?                      �?      �?        颋.���?/�袋.�?      �?        y�5���?�5��P�?              �?      �?      �?/�袋.�?F]t�E�?�������?�������?              �?      �?                      �?�������?�������?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���whG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKㅔh��B�8         �       
             �?�ڰ����?2           ��@              -                    �?��N(��?B           h�@               
       
             �?|�|k6��?2            �U@               	                    �?�����H�?             "@                                  �n@      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �?$��m��?,            �S@                                  T@ZՏ�m|�?            �H@        ������������������������       �                     @                                   �? �#�Ѵ�?            �E@                                   �O@�IєX�?             1@       ������������������������       �                     *@                                   �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                  `X@ ��WV�?             :@        ������������������������       �                     �?        ������������������������       �                     9@               ,                    �?J�8���?             =@                                 �^@�n_Y�K�?             :@                                  �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               )                    �?�X����?             6@              $                   �m@�q�q�?             2@               #                   �a@����X�?             @                      	             �?�q�q�?             @        ������������������������       �                     �?        !       "                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        %       (                    �?�C��2(�?             &@        &       '                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        *       +                     M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        .       c                    �?T�~���?           `{@        /       <                   �f@��N(��?m            �e@        0       9       	          `ff@      �?,             P@       1       8       	          ����?��v$���?*            �N@       2       7                   `X@�?�|�?            �B@        3       4                    �K@r�q��?             @        ������������������������       �                     @        5       6                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ?@        ������������������������       �                     8@        :       ;                     L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        =       L                    �?�{���2�?A            �[@        >       C                   �\@^�!~X�?            �J@        ?       B                    @I@�	j*D�?             *@        @       A                    \@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        D       E                    �?��(\���?             D@        ������������������������       �                     "@        F       G       	          833�?��a�n`�?             ?@        ������������������������       �        	             0@        H       K                   b@z�G�z�?
             .@       I       J       	          ����?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        M       X                   ``@��o	��?#             M@        N       W                   Xp@�q�q�?             8@       O       V                    �I@�����?             5@       P       Q                   �\@r�q��?             (@        ������������������������       �                     �?        R       U                    i@�C��2(�?             &@        S       T       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        Y       Z                    @������?             A@        ������������������������       �                     .@        [       \                   �a@D�n�3�?             3@        ������������������������       �                      @        ]       ^       
             �?���!pc�?             &@        ������������������������       �                     @        _       `                   �d@      �?              @        ������������������������       �                     @        a       b                   p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        d       �                    �P@4�dS���?�            pp@       e       �       	          ����?�U�:��?�            �m@       f       k                   e@�G�V�e�?R             a@        g       h       	          033�?`Ql�R�?             �G@       ������������������������       �                     D@        i       j                    �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        l       q                   �[@NKF����?2            @V@        m       p                    �?���Q��?             $@       n       o       	             �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        r       s                   Pf@p#�����?,            �S@        ������������������������       �                     �?        t                           @N@�ݜ�?+            �S@       u       ~                   �a@�>����?              K@       v       y                    �C@������?            �B@        w       x                    �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        z       }                    \@�#-���?            �A@        {       |                   �`@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     >@        ������������������������       �        
             1@        �       �                    �N@      �?             8@        ������������������������       �                     @        �       �                   p`@ףp=
�?
             4@        �       �                    _@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        �       �                   �W@p���??             Y@        ������������������������       �                     �?        �       �                    �?`�LVXz�?>            �X@       ������������������������       �        .            �R@        �       �                     K@ �q�q�?             8@        �       �       
             �?      �?             @        ������������������������       �                     �?        �       �                   �n@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     ;@        �       �                    �?�=fL�?�            �x@        �       �                    �P@naԵ̗�?S            �`@       �       �                    P@q*� �?O            �_@        �       �                    �M@>���Rp�?             =@       �       �                   �\@���N8�?             5@        �       �                    �?      �?             @       �       �                   `Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        �       �       	          ���@      �?              @       �       �                   �\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?j�Je���?<            �X@        �       �       	          ����?��.k���?             A@       �       �                    �?      �?             8@       �       �                   �q@�q�q�?             5@       �       �                    @F@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        �       �       	          @33�?���Q��?             $@       �       �                   �r@      �?              @        ������������������������       �                     @        �       �                    @M@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �m@�q�q�?             @        ������������������������       �                     �?        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    `P@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?     ��?)             P@       �       �                    �?^�!~X�?"            �J@        ������������������������       �                      @        �       �                    @D@���V��?            �F@        �       �                   �p@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    ]@������?            �D@        �       �                   �k@�	j*D�?             *@        ������������������������       �                     @        �       �                   �[@      �?              @        ������������������������       �                     @        �       �                   �b@z�G�z�?             @       �       �                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        �       �       	          `ff�?�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          033�?��ɉ�?�            @p@       �       �                   �g@���J��?�            �o@       �       �                    c@ ���z��?�            �o@       �       �                   Hp@@9����?�            �l@       ������������������������       �        e             f@        �       �                   @_@���J��?"            �I@        �       �                   �^@�nkK�?             7@       ������������������������       �                     6@        ������������������������       �                     �?        ������������������������       �                     <@        �       �                   Pc@ȵHPS!�?             :@        ������������������������       �                      @        �       �                    �? �q�q�?             8@        �       �                    @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     4@        ������������������������       �                     �?        �       �                    @K@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  �z��A�?����?�>���T�?F0���j�?�2)^ �?;���C��?�q�q�?�q�q�?      �?      �?      �?      �?              �?      �?                      �?              �?�N��N��?vb'vb'�?�>4և��?9/����?              �?�/����?�}A_Ч?�?�?      �?              �?      �?              �?      �?        O��N���?;�;��?              �?      �?        |a���?�rO#,��?ى�؉��?;�;��?      �?      �?              �?      �?        ]t�E]�?�E]t��?UUUUUU�?UUUUUU�?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        F]t�E�?]t�E�?�������?�������?              �?      �?                      �?      �?      �?              �?      �?                      �?�a�]�?��'����?�>���T�?F0���j�?      �?      �?;ڼOqɐ?.�u�y�?к����?*�Y7�"�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?        �9	ą��?,c��2�?�	�[���?�}�	��?;�;��?vb'vb'�?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?�������?              �?�c�1Ƹ?�s�9��?              �?�������?�������?;�;��?�؉�؉�?      �?                      �?      �?        ������?���{�?UUUUUU�?�������?=��<���?�a�a�?�������?UUUUUU�?              �?]t�E�?F]t�E�?      �?      �?      �?                      �?      �?              �?                      �?�?xxxxxx�?              �?(������?l(�����?              �?F]t�E�?t�E]t�?      �?              �?      �?      �?              �?      �?      �?                      �?���w�?*C����?�pR�屵?�A�I�?�������?�������?W�+�ɕ?}g���Q�?              �?�$I�$I�?۶m۶m�?              �?      �?        �9�as�?��g<��?333333�?�������?      �?      �?              �?      �?              �?        �#{���?7a~W��?      �?        �i�i�?\��[���?h/�����?�Kh/��?к����?��g�`��?      �?      �?              �?      �?        _�_�?�A�A�?333333�?�������?              �?      �?                      �?              �?      �?      �?      �?        �������?�������?�$I�$I�?�m۶m��?              �?      �?                      �?{�G�z�?\���(\�?      �?        [�R�֯�?�~�@��?              �?UUUUUU�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?h`Ef��?_~��f��?�}s���?A�d�?�T*�J��?�V��j��?GX�i���?�i��F�?�a�a�?��y��y�?      �?      �?      �?      �?              �?      �?                      �?              �?      �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?x9/���?����>�?�?�������?      �?      �?UUUUUU�?UUUUUU�?]t�E�?F]t�E�?              �?      �?        �������?333333�?      �?      �?              �?�������?333333�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �������?�������?              �?      �?             ��?      �?�}�	��?�	�[���?      �?        [�[��?�>�>��?      �?      �?              �?      �?        �|����?������?vb'vb'�?;�;��?      �?              �?      �?      �?        �������?�������?      �?      �?      �?                      �?              �?      �?        ]t�E�?t�E]t�?      �?                      �?              �??�?��? �����?______�?�?�����~�?�@ �?�}���?p�}�q?      �?        ______�?�?�Mozӛ�?d!Y�B�?      �?                      �?      �?        ��N��N�?�؉�؉�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?�������?333333�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��(hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@>         �                    �?�HK��x�?9           ��@              w                    �?&��f���?;           �@              B       
             �?����?�            �v@                                  �?�TG!u�?�            �n@                      	          `ff�?p9W��S�?             C@                                  @M@r�q��?             8@                                 �a@D�n�3�?             3@              	                   �Z@"pc�
�?             &@        ������������������������       �                     �?        
                          �n@ףp=
�?             $@                      	          ����?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  �b@      �?              @       ������������������������       �                     @                                  `^@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     ,@               A                   �e@�R��ݽ?�             j@              ,                    �?0G���ջ?�             j@               )                    �?�J�4�?              I@                                  �?�Ra����?             F@                                   @P@      �?              @       ������������������������       �                     @                      	          tff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                    @H@�����H�?             B@        ������������������������       �        	             ,@        !       $                   �^@"pc�
�?             6@        "       #                   q@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        %       &                    �K@�r����?	             .@       ������������������������       �                     $@        '       (       	          ����?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        *       +                    @N@      �?             @        ������������������������       �                     @        ������������������������       �                     @        -       >                   0c@pY���D�?e            �c@       .       /       
             �?П��o�?c            `c@        ������������������������       �                     9@        0       1                    `@0�ޤ��?U            @`@        ������������������������       �                    �B@        2       7                   �`@�g�y��?8            @W@        3       6                   �X@���}<S�?             7@        4       5                   l@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             3@        8       9                   pl@`����֜?,            �Q@       ������������������������       �                     E@        :       =                   �[@h�����?             <@        ;       <                   �a@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     2@        ?       @       	             @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        C       J                    �?d%@�"�?D            @]@        D       E                    @M@@4և���?             ,@       ������������������������       �                     $@        F       G                   �p@      �?             @        ������������������������       �                      @        H       I                    e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        K       l                    �?���g�?8            �Y@       L       [       	          ����?z\�3�?*            �S@       M       T                    �?@�r-��?            �M@        N       S                   f@�z�G��?             4@        O       R                    �L@      �?              @       P       Q                   �[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        U       Z                   �e@$�q-�?            �C@       V       W                   �c@�?�|�?            �B@       ������������������������       �                     >@        X       Y                     H@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        \       e                     L@�G�z��?             4@       ]       ^                   0`@�q�q�?             (@        ������������������������       �                      @        _       `                    �?�z�G��?             $@        ������������������������       �                     �?        a       d                   0l@�<ݚ�?             "@        b       c                    �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        f       g       	            �?      �?              @        ������������������������       �                      @        h       i                    �?�q�q�?             @        ������������������������       �                     �?        j       k                   �]@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        m       v                   pf@r�q��?             8@       n       o                    �?�C��2(�?             6@       ������������������������       �                     0@        p       u                     P@�q�q�?             @       q       r                   �`@�q�q�?             @        ������������������������       �                     �?        s       t                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        x       �                    �?��<�Ұ?X            `b@       y       �                    `R@��ɹ?;            �W@       z       �                    �?H��2�?:            @W@        {       �       	          833�? >�֕�?            �A@        |       }                   0`@"pc�
�?             &@       ������������������������       �                     @        ~                          �c@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     8@        �       �                   �p@XB���?%             M@       ������������������������       �                     I@        �       �                   `@      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �J@        �       �                   �b@���և�?�            py@       �       �       
             �?Z�U��?�             k@        �       �       	          ���@�s�n_�?>             Z@       �       �                    �?�C+����?=            @Y@        �       �                     P@�\��N��?             3@       �       �                    �I@�	j*D�?             *@        ������������������������       �                     @        �       �                   @]@���Q��?             $@        �       �                   �u@r�q��?             @       �       �                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �n@�p ��?2            �T@       �       �                    �?�<ݚ�?&             K@        �       �                   �^@և���X�?             @        �       �                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �X@t/*�?!            �G@        �       �                   �W@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �c@,���i�?            �D@       �       �                   �`@�˹�m��?             C@       ������������������������       �                     6@        �       �                   �m@     ��?             0@       �       �                   �\@�r����?             .@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        �       �                    �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     <@        ������������������������       �                     @        �       �                    @L@ d�=��?G            @\@       �       �       	          ����?�|���?7             V@       ������������������������       �        3             T@        �       �                    g@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    p@ �o_��?             9@       �       �                    �Q@      �?
             0@       ������������������������       �                     ,@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @Q@�q�q�?             "@       �       �                     @؇���X�?             @        �       �                   0b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�?�'�@�?y            �g@        �       �       
             �?      �?&             P@        �       �                    �?      �?             0@       �       �                   �g@z�G�z�?
             .@        �       �                    @G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     H@        �       �                    �F@r�q��?S            �_@        �       �                    d@h㱪��?#            �K@        �       �                    @�<ݚ�?             "@       �       �                   Hp@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     G@        �       �                   �e@���BK�?0            �Q@       �       �                   �t@�J�4�?#             I@       �       �                   �n@؇���X�?"            �H@       �       �                   �l@��a�n`�?             ?@       �       �                    @M@HP�s��?             9@       ������������������������       �                     2@        �       �                    j@����X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �m@r�q��?             @       ������������������������       �                     @        �       �                   0n@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        �       �       
             �?�G��l��?             5@        �       �                   @b@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �                    f@���|���?	             &@       �       �                    �L@�<ݚ�?             "@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �T8q���?��cG��?ҤI�&M�?˖-[�l�?R�Q��?Ws5Ws5�?�����߸?@�O%��?l(�����?�k(����?UUUUUU�?UUUUUU�?l(�����?(������?/�袋.�?F]t�E�?              �?�������?�������?�������?�������?              �?      �?              �?              �?      �?              �?      �?      �?              �?      �?                      �?              �?ϧ��د?��#s�?�؉�؉�?vb'vb'�?{�G�z�?�z�G��?]t�E�?]t�E]�?      �?      �?              �?      �?      �?      �?                      �?�q�q�?�q�q�?              �?F]t�E�?/�袋.�?�$I�$I�?�m۶m��?              �?      �?        �?�������?              �?�������?333333�?              �?      �?              �?      �?              �?      �?        �3���?a~W��0�?�=�ѓ?a�qa�?              �?z�z��?/�B/�B�?              �?�B!��?��{���?d!Y�B�?ӛ���7�?      �?      �?      �?                      �?              �?�A�A�?�������?              �?�$I�$I�?�m۶m��?�������?�������?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �LɔL��?�fm�fm�?n۶m۶�?�$I�$I�?      �?              �?      �?      �?              �?      �?              �?      �?        ^�	���?C����?��jq��?h *�3�?'u_�?��c+���?ffffff�?333333�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        �؉�؉�?;�;��?*�Y7�"�?к����?      �?        ۶m۶m�?�$I�$I�?      �?                      �?              �?�������?�������?�������?�������?              �?ffffff�?333333�?              �?9��8���?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?        UUUUUU�?�������?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?        [��5;j�?�7�L\��?m�w6�;�?���\AL�?X`��?�~�駟�?�A�A�?��+��+�?F]t�E�?/�袋.�?              �?      �?      �?      �?                      �?              �?�{a���?GX�i���?              �?      �?      �?      �?                      �?      �?                      �?�6��1�?'������?��LW�+�?͢fQ���?O��N���?��N��N�?��g����?&���?y�5���?�5��P�?;�;��?vb'vb'�?              �?�������?333333�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?      �?                      �?      �?        ��+Q��?Q��+Q�?�q�q�?9��8���?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        W�+���?�;����?      �?      �?              �?      �?        8��18�?�����?^Cy�5�?��P^Cy�?              �?      �?      �?�?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ���	��?x�!���?��.���?F]t�E�?      �?              �?      �?              �?      �?        
ףp=
�?�Q����?      �?      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        ������?y�5���?      �?      �?      �?      �?�������?�������?      �?      �?      �?                      �?      �?                      �?      �?        �������?UUUUUU�?־a���?��)A��?9��8���?�q�q�?      �?      �?      �?                      �?              �?      �?        ��RO�o�?$Zas �?�z�G��?{�G�z�?۶m۶m�?�$I�$I�?�c�1��?�s�9��?q=
ףp�?{�G�z�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?                      �?��y��y�?1�0��?333333�?ffffff�?              �?      �?        ]t�E]�?F]t�E�?9��8���?�q�q�?      �?      �?      �?                      �?              �?              �?�t�bub��)     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���PhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         �                    �?�7i���?U           ��@              q       	          `ff�?<�_����?�           ��@              0       
             �?�O:���?           �z@                                  �c@�z��W�?K            �\@        ������������������������       �                    �@@                                   �?^�JB=�?7            @T@               
                   `m@�n_Y�K�?             :@               	                    @N@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @                                   _@��.k���?             1@        ������������������������       �                     @                      	            �?և���X�?
             ,@                                  �?�q�q�?	             (@                                 pb@      �?              @        ������������������������       �                     @                                   �J@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @               )                    �O@���!pc�?%            �K@              (                   (q@���V��?            �F@              !                   �b@     ��?             @@                                 �a@���7�?             6@       ������������������������       �                     1@                      	          ����?z�G�z�?             @        ������������������������       �                     @                                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        "       '                   0a@���Q��?             $@       #       $                   0e@      �?              @       ������������������������       �                     @        %       &                   �f@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        *       /                    �P@z�G�z�?             $@       +       ,                    �?�����H�?             "@       ������������������������       �                     @        -       .                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        1       H                    �?lΜT ��?�            ps@        2       E       	          ����?~���L0�?"            �H@       3       B                   �q@���y4F�?             C@       4       5                    `@ףp=
�?             >@        ������������������������       �                     @        6       ?       	          ����?�LQ�1	�?             7@       7       >                    m@�����?             5@        8       =                    @L@      �?              @       9       <                   i@؇���X�?             @        :       ;                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             *@        @       A                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        C       D                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        F       G                   pb@���|���?             &@       ������������������������       �                     @        ������������������������       �                     @        I       T                    I@��L�$�?�            `p@        J       M                    ^@���Q��?             .@        K       L                   @U@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        N       O                    �?X�<ݚ�?             "@        ������������������������       �                     @        P       S                   �b@r�q��?             @       Q       R                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        U       f                    �?М�x�2�?�            �n@        V       e                    �?h�WH��?%             K@       W       ^                    b@,���i�?            �D@       X       Y                    �?�IєX�?             A@       ������������������������       �                     <@        Z       ]                    a@�q�q�?             @       [       \                    @K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        _       `                    j@և���X�?             @        ������������������������       �                      @        a       b                    �?z�G�z�?             @        ������������������������       �                     �?        c       d                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        g       h                    @L@@��A� �?w             h@       ������������������������       �        h             e@        i       j                   `a@�8��8��?             8@        ������������������������       �                     (@        k       l                    �?r�q��?	             (@        ������������������������       �                     @        m       n                   0b@����X�?             @        ������������������������       �                     �?        o       p                    �N@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        r       �       
             �?4�c���?�            �r@       s       �                    �?�L����?�            @o@        t       �       	          `ff�?��Q:��?*            �M@       u       �       	          ����?f���M�?             ?@       v       w                    @F@�eP*L��?             6@        ������������������������       �                     @        x       }                    �K@j���� �?             1@        y       z                   �^@      �?              @        ������������������������       �                     @        {       |                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ~                          �W@�q�q�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                   �`@���Q��?             @        ������������������������       �                      @        �       �                   xu@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�����H�?             "@        �       �                   `]@�q�q�?             @        ������������������������       �                     �?        �       �                    @P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �l@@4և���?             <@        �       �                    �?z�G�z�?             $@        �       �                   0`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        �       �                    �?�g$����?{            �g@       �       �       	          ����?�7��?e            �c@        �       �                   �`@�GN�z�?             6@       �       �                    @L@     ��?             0@       �       �                   �r@������?
             .@       �       �                    @G@r�q��?             (@       �       �                   �j@�q�q�?             @        ������������������������       �                      @        �       �                   @n@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Z@��J��i�?U            �`@        ������������������������       �                     �?        �       �       	          `ff @���%yU�?T            �`@       �       �                    @M@pY���D�?2            �S@       ������������������������       �        $            �M@        �       �                   �p@ףp=
�?             4@       ������������������������       �        
             ,@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        "             K@        �       �                   P`@">�֕�?            �A@        �       �                    �?���Q��?
             .@        ������������������������       �                     @        �       �                   �\@      �?	             (@        ������������������������       �                      @        �       �                   `_@���Q��?             $@        ������������������������       �                     @        �       �       	             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �T@ףp=
�?             4@        �       �                   �d@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     *@        �       �       	          ���@�J��%�?            �H@       �       �                    �?������?            �F@       �       �                    c@և���X�?             5@       �       �                    �H@�t����?             1@        �       �                   ph@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    S@8�Z$���?             *@        �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�C��2(�?	             &@        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                     @        �       �                   p`@��3��?            @h@        �       �                    �?ą%�E�?9            @V@       �       �       
             �?��?^�k�?.            �Q@       ������������������������       �        "            �J@        �       �                    �?�t����?             1@       �       �                    ]@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                   �Y@p�ݯ��?             3@        ������������������������       �                      @        �       �                   @_@���|���?             &@       ������������������������       �                     @        �       �                   �c@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �I@�n����?F            @Z@        �       �                    �?�	j*D�?             *@        ������������������������       �                      @        �       �                    �?"pc�
�?             &@       �       �                    @G@      �?              @        ������������������������       �                     @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?��H�?>             W@       �       �                   �a@XB���?&             M@        �       �                   �u@�C��2(�?             6@       ������������������������       �                     4@        ������������������������       �                      @        ������������������������       �                     B@        �       �       	          ����?�ʻ����?             A@       �       �       
             �?      �?             4@        �       �       	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             (@        ������������������������       �        
             ,@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  }}}}}}�?AAAAAA�?�<�0&�?]��ҟ��?��
>q��?�P���?u�YLg�?�t�YL�?              �?�2�tk~�?��E���?;�;��?ى�؉��?9��8���?�q�q�?      �?                      �?�������?�?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?      �?              �?333333�?�������?      �?                      �?      �?      �?      �?                      �?      �?        t�E]t�?F]t�E�?�>�>��?[�[��?      �?      �?F]t�E�?�.�袋�?              �?�������?�������?              �?      �?      �?      �?                      �?333333�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�������?�������?�q�q�?�q�q�?      �?              �?      �?      �?                      �?              �?��0�t�?y{�X�?����>4�?������?6��P^C�?(������?�������?�������?      �?        ��Moz��?Y�B��?=��<���?�a�a�?      �?      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?      �?              �?      �?              �?      �?              �?      �?        F]t�E�?]t�E]�?              �?      �?        �:�ֆi�?�U���g�?333333�?�������?�������?UUUUUU�?              �?      �?        �q�q�?r�q��?      �?        UUUUUU�?�������?      �?      �?              �?      �?                      �?}����?S���.�?��^B{	�?B{	�%��?�����?8��18�?�?�?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?              �?      �?              �?      �?              �?        �/����?��H	9�?      �?        UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?6�TWέ�?3�*j��?ˡE����?��n���?�A�I��?'u_[�?��RJ)��?��Zk���?t�E]t�?]t�E�?      �?        ZZZZZZ�?�������?      �?      �?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?        �$I�$I�?n۶m۶�?�������?�������?      �?      �?      �?                      �?      �?      �?      �?                      �?              �?T��Iw�?���?�A�A�?��[��[�?]t�E�?�袋.��?      �?      �?�?wwwwww�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?���@��?�[�՘H�?      �?        ���̎?M�3�τ�?�3���?a~W��0�?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�A�A�?_�_��?333333�?�������?      �?              �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�$I�$I�?�m۶m��?              �?      �?                      �?c}h���?9/����?wwwwww�?�?۶m۶m�?�$I�$I�?�������?�������?      �?      �?      �?                      �?;�;��?;�;��?      �?      �?              �?      �?        F]t�E�?]t�E�?      �?      �?      �?                      �?              �?      �?              �?                      �?W?���?*���:�?��g<�?�as���?�A�A�?_�_��?              �?�?<<<<<<�?�$I�$I�?�m۶m��?              �?      �?                      �?Cy�5��?^Cy�5�?              �?]t�E]�?F]t�E�?      �?        �������?�������?              �?      �?         �����?8�8��?vb'vb'�?;�;��?              �?/�袋.�?F]t�E�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        zӛ����?!Y�B�?�{a���?GX�i���?F]t�E�?]t�E�?              �?      �?                      �?<<<<<<�?�������?      �?      �?      �?      �?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ@f�"hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�>         B                   �_@�>���?/           ��@                      	            �?�r&��K�?w            `g@                                   �?�1��u�?0            @R@                                 �e@d}h���?#             L@              
                    �?z�G�z�?"            �K@                     
             �?@-�_ .�?            �B@       ������������������������       �                     A@               	       	          `ffֿ�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   @      �?
             2@                                  U@      �?             (@        ������������������������       �                      @                                   �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                   [@��.k���?             1@        ������������������������       �                     @                                   �P@�n_Y�K�?	             *@                                  �?���!pc�?             &@                                  �?z�G�z�?             $@        ������������������������       �                     @                                  �\@      �?             @        ������������������������       �                     �?                                   a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                ?                   �c@l�b�G��?G            �\@       !       6                    �? ѯ��?C            �Z@       "       +       
             �?`��F:u�?7            �U@       #       *                   �_@P����?'            �M@        $       )                    �?P���Q�?             4@        %       (       	             �?�����H�?             "@       &       '                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                    �C@        ,       -       	          033�? �Cc}�?             <@        ������������������������       �                     "@        .       3                    �?�S����?
             3@       /       0                     M@��S�ۿ?             .@        ������������������������       �                     @        1       2                    @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        4       5                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        7       8                   @_@ףp=
�?             4@        ������������������������       �                     $@        9       :       
             �?z�G�z�?             $@        ������������������������       �                     �?        ;       <                    �?�����H�?             "@        ������������������������       �                      @        =       >                    ]@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        @       A       	          033@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        C       �                    �?pxE'��?�           ؆@       D       s                    �?��w(���?           �}@        E       `       	          pff�?և���X�?U            `b@       F       M       
             �?�j<,���?=            @[@        G       H       	          ����?RB)��.�?            �E@       ������������������������       �                     @@        I       J                   �p@"pc�
�?             &@       ������������������������       �                     @        K       L                   �c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        N       Y                    �L@���!pc�?$            �P@       O       R                   `i@�LQ�1	�?             G@        P       Q                    ^@      �?              @        ������������������������       �                     @        ������������������������       �                     @        S       X                    �?P�Lt�<�?             C@       T       W                    l@ 7���B�?             ;@        U       V                    a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     8@        ������������������������       �                     &@        Z       [                   �b@���Q��?
             4@        ������������������������       �                     @        \       ]                   @d@$�q-�?             *@        ������������������������       �                     @        ^       _                    _@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        a       l                    �N@�S����?             C@       b       k                    �?ܷ��?��?             =@       c       d                    �?��2(&�?             6@        ������������������������       �                     @        e       j       
             �?     ��?             0@       f       g                   hq@@4և���?
             ,@       ������������������������       �                     $@        h       i                    �J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        m       r                     P@�q�q�?             "@       n       q                    �?���Q��?             @       o       p                   �q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        t       �       	          033�?���O1��?�            �t@       u       v                   �W@`�^�
�?�            s@        ������������������������       �                     @        w       �       
             �?(+ �8�?�            �r@        x       �                    �?��y�:�?(            �P@       y       �       	          ����?z�G�z�?"            �K@        z       {                   @b@      �?
             ,@        ������������������������       �                     @        |       }                   �n@�z�G��?             $@        ������������������������       �                     @        ~                           _@���Q��?             @        ������������������������       �                      @        �       �                   8p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?������?            �D@        �       �                   �^@�θ�?             *@        �       �                     I@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?h�����?             <@       ������������������������       �                     6@        �       �                    �M@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�8��8��?             (@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                    @�/�!�?�            `m@       �       �       	            �?�HGݐ\�?�            `k@       ������������������������       �        m             f@        �       �                   �_@�����?             E@        �       �                    �D@և���X�?             @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �A@        �       �                   ``@     ��?             0@        �       �                    ^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                   �`@�5��?             ;@       �       �                    �L@     ��?             0@       �       �                   �^@      �?	             (@        �       �                    c@���Q��?             @       �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        �       �       
             �?�9���[�?�            �o@       �       �                   P`@��JB��?�            �i@        �       �       	          ����?�������?1             V@       �       �                    @L@     ��?!             P@       �       �                    �?<���D�?            �@@        �       �                   @_@      �?             @        ������������������������       �                      @        �       �       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          ����?XB���?             =@       ������������������������       �                     8@        �       �                   m@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?`՟�G��?             ?@        �       �       	             �?      �?              @       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ]@\X��t�?             7@        ������������������������       �                     @        �       �       	          ����?      �?
             4@       �       �                   �[@�q�q�?             .@        ������������������������       �                     @        �       �                   `]@      �?             $@        ������������������������       �                     @        �       �       	             �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@        �       �       	          ����?T(y2��?P            �]@        �       �                   �n@�������?             >@        �       �                    �K@�eP*L��?	             &@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   ``@r�q��?             @       ������������������������       �                     @        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�KM�]�?             3@        �       �       	          ����?�<ݚ�?             "@        �       �                    d@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                   `c@ }�Я��?:            @V@       ������������������������       �        9             V@        ������������������������       �                     �?        �       �       	          ����?��S���?            �F@       �       �                   `@r֛w���?             ?@        ������������������������       �                     (@        �       �                   �n@D�n�3�?             3@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���|���?             &@       �       �                    �?      �?              @       ������������������������       �                     @        �       �                   @d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?@4և���?	             ,@       �       �                   �p@ףp=
�?             $@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �Kh/��?��Kh/�?*�Ap*�?5{��c5�?�1bĈ�?�s�Ν;�?۶m۶m�?I�$I�$�?�������?�������?к����?S�n0E�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?�������?�������?      �?                      �?              �?      �?        �?�������?              �?;�;��?ى�؉��?F]t�E�?t�E]t�?�������?�������?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?p�}��?�Gp��?�@�Ե�?n���4�?Ȥx�L��?�u�7[��?'u_[�?�V'u�?�������?ffffff�?�q�q�?�q�q�?�������?�������?              �?      �?                      �?              �?              �?۶m۶m�?%I�$I��?              �?^Cy�5�?(������?�?�������?              �?      �?      �?      �?                      �?      �?      �?      �?                      �?�������?�������?              �?�������?�������?      �?        �q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?      �?                      �?�$I�$I�?�m۶m��?              �?      �?        I=C�a�?n�y�=�?̾�2.�?h�t���?۶m۶m�?�$I�$I�?����?���]8��?���)k��?S֔5eM�?              �?/�袋.�?F]t�E�?      �?              �?      �?      �?                      �?F]t�E�?t�E]t�?��Moz��?Y�B��?      �?      �?              �?      �?        ���k(�?(�����?	�%����?h/�����?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?        �������?333333�?      �?        ;�;��?�؉�؉�?              �?�$I�$I�?۶m۶m�?      �?                      �?^Cy�5�?(������?a���{�?��=���?t�E]t�?��.���?              �?      �?      �?�$I�$I�?n۶m۶�?              �?      �?      �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?333333�?�������?      �?      �?              �?      �?                      �?              �?P�M�_�?���ˊ��?�m����?^���ۺ?              �?g���Y��?�Tb*1��?�@��~�?~5&��?�������?�������?      �?      �?              �?ffffff�?333333�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        �|����?������?ى�؉��?�؉�؉�?�������?333333�?      �?                      �?      �?        �m۶m��?�$I�$I�?      �?        �������?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?�]~���?J4p���?����_j�?@+���?      �?        =��<���?�a�a�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?�������?333333�?              �?      �?              �?              �?      �?      �?      �?      �?                      �?      �?        /�����?h/�����?      �?      �?      �?      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?F]t�E�?/�袋.�?      �?                      �?Y�eY�e�?j��i���?�{����?ᖚ��?/�袋.�?t�E]t�?      �?      �?|���?|���?      �?      �?      �?              �?      �?              �?      �?        �{a���?GX�i���?              �?�������?�������?      �?                      �?�s�9��?�1�c��?      �?      �?      �?      �?              �?      �?                      �?!Y�B�?��Moz��?      �?              �?      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?�������?UUUUUU�?              �?      �?                      �?              �?�5�5�?�F��F��?�������?�������?]t�E�?t�E]t�?�������?�������?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?(�����?�k(���?�q�q�?9��8���?      �?      �?              �?      �?                      �?              �?p�\��?�я~���?              �?      �?        �?�������?���{��?�B!��?      �?        l(�����?(������?      �?      �?              �?      �?        F]t�E�?]t�E]�?      �?      �?              �?      �?      �?              �?      �?              �?        �$I�$I�?n۶m۶�?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��O,hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKㅔh��B�8         r                    �?�LT ���?9           ��@                                  �B@�%�Gt@�?2           �~@                                   �?������?             .@                                 `]@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @               9       	          033�?���c��?,           �}@        	       
                   �X@�û��|�?x             g@        ������������������������       �                     4@                       
             �?�>$�*��?m            �d@                                  @J@P�;�&��?9            @U@                      	          833�?@-�_ .�?            �B@       ������������������������       �                     =@                                   �?      �?              @        ������������������������       �                      @        ������������������������       �                     @                                  @l@      �?              H@                                  b@XB���?             =@       ������������������������       �                     8@                                  �_@z�G�z�?             @        ������������������������       �                      @                                  �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                      	          ����?D�n�3�?             3@        ������������������������       �                     @                                  �]@8�Z$���?             *@                                  �[@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        !       ,                   �b@ܩ�d	��?4            �S@       "       #                   `\@��ϭ�*�?%             M@        ������������������������       �        	             1@        $       +       	          ����?,���i�?            �D@       %       &                    �?�?�|�?            �B@       ������������������������       �                    �@@        '       (                    �?      �?             @        ������������������������       �                      @        )       *       	          833�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        -       0                    �?���N8�?             5@        .       /                    @M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        1       8                    �K@�t����?             1@       2       7                   �f@"pc�
�?             &@       3       6                   �[@ףp=
�?             $@        4       5                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        :       S       	          ����?�B#�{�?�            @r@        ;       J                    �?�+$�jP�?2            @T@       <       C                   �c@X��Oԣ�?%             O@       =       B                   �[@ 7���B�?!             K@        >       ?                    �H@����X�?             @        ������������������������       �                     @        @       A                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �G@        D       I                    �?      �?              @       E       H                   �`@����X�?             @       F       G                   �e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        K       L                   �i@D�n�3�?             3@       ������������������������       �                     "@        M       R                   �q@z�G�z�?             $@       N       O                    ^@���Q��?             @        ������������������������       �                      @        P       Q                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        T       k                   @e@0�ڂcv�?�            `j@       U       h                    �R@��)Cd�?~            �i@       V       a                   �_@P����֨?|             i@        W       \                   �^@ ,��-�?!            �M@       X       Y       
             �?@3����?             K@       ������������������������       �                     I@        Z       [       	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ]       `                   0p@���Q��?             @       ^       _                    �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        b       c                   q@ ��U��?[            �a@       ������������������������       �        =            �W@        d       e                     M@@��8��?             H@       ������������������������       �                     7@        f       g                   Xq@`2U0*��?             9@        ������������������������       �                     �?        ������������������������       �                     8@        i       j                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        l       m                    �?���Q��?             @        ������������������������       �                      @        n       q                    �?�q�q�?             @       o       p       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        s       �                   �`@�*�g`�?           �z@        t       �                   @c@
XU�)��?M            �_@        u       �                    `@�q��/��?            �H@       v       �                    �?�����?             E@        w       �       	          033�?z�G�z�?             4@       x       �                    ^@      �?	             0@       y       �                    �O@����X�?             @       z       {       	             �r�q��?             @        ������������������������       �                     �?        |                           �?z�G�z�?             @       }       ~                    \@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �       
             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        �       �                   `_@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?$��m��?1            �S@        �       �                    �?V������?            �B@        ������������������������       �                     $@        �       �                    �? 7���B�?             ;@        �       �                    @M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     8@        �       �                    �?��Y��]�?            �D@       ������������������������       �                    �A@        �       �                     P@r�q��?             @        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @L@j�q����?�            �r@       �       �                   �c@�^����?�            �m@        �       �       	          ����?�n_Y�K�?             *@       �       �                     B@z�G�z�?             $@        �       �                     @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          033�?@�@+��?�            �k@       �       �       	          ����?��qn�H�?            �i@       �       �                    �?�h����?k             e@       �       �                   @g@`���i��?;             V@       ������������������������       �        :            �U@        ������������������������       �                      @        �       �                    @E@p=
ףp�?0             T@        ������������������������       �                     C@        �       �                   �q@r�q��?             E@       �       �       	          ����?�KM�]�?             C@       �       �                    �?؇���X�?             <@       �       �                    �H@�����H�?             ;@        �       �       
             �?      �?             (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �        	             .@        ������������������������       �                     �?        ������������������������       �        	             $@        �       �                   �r@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �d@�S����?             C@       �       �                   �b@     ��?             @@       �       �                   0a@(;L]n�?             >@       ������������������������       �                     ;@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ^@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?��.k���?
             1@       �       �                   `d@�q�q�?             (@        ������������������������       �                     @        �       �                    @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    a@     ��?*             P@        �       �                   �r@�q�q�?             5@       �       �       	          ����?�<ݚ�?             2@        �       �                    `@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    `@�C��2(�?             &@       ������������������������       �                     @        �       �                   @c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �P@^����?            �E@       �       �       	          ����?���@��?            �B@        �       �                   �b@��.k���?             1@       �       �                    d@      �?	             (@       �       �                     P@      �?              @       �       �                    @N@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B0  ��u���?�(E~��?ئ@���?J���?wwwwww�?�?;�;��?;�;��?              �?      �?                      �?{1�z1��?�3X�3X�?��,d!�?8��Moz�?              �?�����?�18���?�?�������?к����?S�n0E�?              �?      �?      �?      �?                      �?      �?      �?�{a���?GX�i���?              �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?l(�����?(������?              �?;�;��?;�;��?333333�?�������?      �?                      �?      �?        ��7a~�?�ґ=�?����=�?|a���?      �?        �����?8��18�?*�Y7�"�?к����?      �?              �?      �?      �?              �?      �?              �?      �?                      �?��y��y�?�a�a�?      �?      �?      �?                      �?�?<<<<<<�?F]t�E�?/�袋.�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�z��ի�?�P�B�
�?B{	�%��?/�����?�s�9�?c�1�c�?h/�����?	�%����?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?      �?      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?(������?l(�����?              �?�������?�������?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �
��T�?Q/#�.�?#>�Tr^�?����?�C��x�?�e0
84�?'u_[�?[4���?h/�����?���Kh�?              �?      �?      �?              �?      �?        333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        ��V�|?���RO��?              �?UUUUUU�?UUUUUU�?              �?{�G�z�?���Q��?      �?                      �?�������?�������?              �?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?{� ���?
����?.���r��?i4�F��?և���X�?/����?�a�a�?=��<���?�������?�������?      �?      �?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?�������?�������?      �?      �?              �?      �?                      �?      �?                      �?      �?      �?              �?      �?                      �?�$I�$I�?�m۶m��?              �?      �?        �N��N��?vb'vb'�?o0E>��?�g�`�|�?      �?        h/�����?	�%����?UUUUUU�?UUUUUU�?              �?      �?                      �?8��18�?������?      �?        �������?UUUUUU�?      �?              �?      �?      �?                      �?=
ףp=�?
ףp=
�?u_[4�?W'u_�?;�;��?ى�؉��?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?������?;Ӹ�Qg�?24��~��?r^�	��?�$I�$I�?۶m۶m�?F]t�E�?F]t�E�?      �?                      �?333333�?ffffff�?      �?        �������?UUUUUU�?�k(���?(�����?۶m۶m�?�$I�$I�?�q�q�?�q�q�?      �?      �?              �?      �?              �?                      �?      �?              �?      �?              �?      �?        (������?^Cy�5�?      �?      �?�������?�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?      �?        �������?�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?�q�q�?9��8���?۶m۶m�?�$I�$I�?      �?                      �?F]t�E�?]t�E�?              �?      �?      �?      �?                      �?      �?        �qG��?w�qG��?L�Ϻ��?к����?�������?�?      �?      �?      �?      �?�������?333333�?      �?                      �?      �?              �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJlBg1hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B�@         (                   p`@SH7�j�?:           ��@                                   @O@��E�"�?o            �f@                     
             �?X�.�d�?U            �a@                                 �X@�ջ����?>             Z@               
                    �?      �?
             0@                                   �?؇���X�?             @       ������������������������       �                     @               	                    V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        4             V@                                  @E@�KM�]�?             C@                                 @b@�X�<ݺ?             B@                     	          ����г�wY;�?             A@        ������������������������       �                     �?        ������������������������       �                    �@@                                   ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                  �`@R���Q�?             D@                                   ^@������?	             .@       ������������������������       �                     $@                                  0`@z�G�z�?             @                                   �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               %                    �Q@HP�s��?             9@                      	          033�?�nkK�?             7@        ������������������������       �                     $@        !       "       
             �?$�q-�?
             *@       ������������������������       �                      @        #       $                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        &       '       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        )       �                    �?�b��f��?�            �@       *       �       	          pff�?ޔ��?           �}@       +       V                    @L@b�?ilX�?�            �w@       ,       9       
             �?P��S�I�?�             q@        -       .                    �?�LQ�1	�?             G@        ������������������������       �                     @        /       8                   �^@      �?             D@       0       1                   �a@�eP*L��?             6@        ������������������������       �                     @        2       3                    �D@�q�q�?	             .@        ������������������������       �                     @        4       7                    �?�C��2(�?             &@        5       6                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        :       O       	          pff�?�Ȍ���?�            �l@       ;       H                   �[@�Ń��̧?�            @j@        <       A                    �?�r����?             >@        =       >                    b@�q�q�?             @        ������������������������       �                      @        ?       @                   �g@      �?             @        ������������������������       �                      @        ������������������������       �                      @        B       C                    �?�8��8��?             8@       ������������������������       �        	             .@        D       G                    �G@�<ݚ�?             "@        E       F                   @[@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        I       J                   �f@ Y@��?m            �f@       ������������������������       �        c            �d@        K       N                    �?      �?
             0@        L       M                   �f@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        P       Q                    �?�q�q�?
             2@        ������������������������       �                     @        R       U                    �J@�eP*L��?             &@       S       T                   0`@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        W       j       
             �?(�-~ ��??            @[@        X       ]                    �?D�n�3�?             C@        Y       \       	          @33�?�����H�?             "@        Z       [                   p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ^       i                   pr@�c�Α�?             =@       _       d                   �a@�J�4�?             9@        `       a                    a@      �?              @        ������������������������       �                     @        b       c                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        e       f                     Q@�IєX�?	             1@       ������������������������       �                     ,@        g       h                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        k       z                    �?�ګH9�?)            �Q@        l       y                    �?j���� �?             1@       m       x                   �b@�q�q�?             (@       n       w       	          ����?X�<ݚ�?             "@       o       r                   �_@      �?              @        p       q                   o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       t                   �d@z�G�z�?             @        ������������������������       �                     @        u       v                   �r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        {       �                   �l@�{��?��?             K@        |       }                    d@���N8�?             5@       ������������������������       �                     0@        ~                           @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �L@:ɨ��?            �@@        �       �                   �`@r�q��?             @        ������������������������       �                     @        �       �                   �n@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     P@�+$�jP�?             ;@       �       �                    d@�q�q�?	             .@       �       �                   �b@      �?             $@       �       �                    @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �       �                   �r@�q�Q�?6             X@       �       �                    �E@��]�T��?-            �T@        �       �                   @a@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �       
             �?����X�?'            �Q@       �       �                    �?z�G�z�?            �K@        ������������������������       �                     7@        �       �                   �a@     ��?             @@       �       �                    �?������?             ;@        �       �       	          033�?����X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       	          `ff�?ףp=
�?             4@       �       �                    �P@z�G�z�?             $@       �       �                   `a@�����H�?             "@       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    @J@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   0b@���Q��?	             .@        �       �                   �n@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    e@      �?              @       ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ���@d}h���?	             ,@       ������������������������       �                     &@        ������������������������       �                     @        �       �       	          033�?�qu�C��?�            p@        �       �                   �b@�ݜ����?#            �M@       �       �                    `@4�B��?            �B@       �       �       	          pff�?      �?             8@       �       �       
             �?�eP*L��?             6@       �       �                   �[@؇���X�?
             ,@        �       �                   �`@�q�q�?             @       ������������������������       �                     @        �       �                   m@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     *@        �       �                    @M@��2(&�?             6@       �       �                    �?�X�<ݺ?             2@        �       �       
             �?      �?              @        ������������������������       �                     @        �       �                   @d@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �j@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   `\@�FVQ&�?�            �h@        �       �       	          033@@�0�!��?             1@       �       �                     M@�r����?             .@       �       �                    b@����X�?             @       �       �                   Pk@      �?             @        ������������������������       �                     �?        �       �                   �m@�q�q�?             @        ������������������������       �                     �?        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �J@PÅ�R1�?}            �f@        �       �                   �c@\-��p�?(             M@       �       �                    �G@�����H�?$             K@        ������������������������       �                     4@        �       �                    `@@�0�!��?             A@       �       �                    �?�����?             5@        �       �                   @[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �_@�}�+r��?             3@        �       �                   �Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     1@        �       �                    b@�	j*D�?             *@       �       �                   �`@ףp=
�?             $@       �       �                   �a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �       	          033@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �? �|ك�?U            �^@       ������������������������       �        N            �[@        �                         `_@�8��8��?             (@        �             	          @33�?�q�q�?             @       �                          �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �t�b�!5     h�h)h,K ��h.��R�(KMKK��hb�B0  ���t��?�~�E)�?����?���?�@�6�?�ۥ����?;�;��?;�;��?      �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?              �?(�����?�k(���?�q�q�?��8��8�?�?�?      �?                      �?      �?      �?      �?                      �?      �?        333333�?333333�?�?wwwwww�?              �?�������?�������?      �?      �?      �?                      �?      �?        {�G�z�?q=
ףp�?d!Y�B�?�Mozӛ�?              �?;�;��?�؉�؉�?              �?�������?�������?      �?                      �?      �?      �?      �?                      �?-d!Y��?�7��Mo�?�!_r��?��A�+�?ǩ��|;�?�X�?t2}�06�?16�='�?d!Y�B�?Nozӛ��?      �?              �?      �?]t�E�?t�E]t�?              �?UUUUUU�?UUUUUU�?              �?]t�E�?F]t�E�?�������?�������?              �?      �?              �?                      �?Lg1��t�?:��,���?��<��<�?�a�a�?�������?�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?        9��8���?�q�q�?      �?      �?              �?      �?              �?        (}�'}��?l�l�v?      �?              �?      �?�������?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?        ]t�E�?t�E]t�?�$I�$I�?۶m۶m�?              �?      �?              �?        D���A�?�w� z|�?(������?l(�����?�q�q�?�q�q�?      �?      �?              �?      �?              �?        �{a���?5�rO#,�?{�G�z�?�z�G��?      �?      �?              �?      �?      �?              �?      �?        �?�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        e�v�'��?6��9�?�������?ZZZZZZ�?�������?�������?r�q��?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?              �?      �?      �?                      �?              �?              �?      �?        ���^B{�?/�����?��y��y�?�a�a�?      �?        �������?�������?      �?                      �?N6�d�M�?e�M6�d�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        /�����?B{	�%��?UUUUUU�?UUUUUU�?      �?      �?�������?UUUUUU�?      �?                      �?              �?      �?              �?        UUUUUU�?UUUUUU�?jW�v%j�?KԮD�J�?�������?UUUUUU�?              �?      �?        �$I�$I�?�m۶m��?�������?�������?              �?      �?      �?{	�%���?B{	�%��?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?�������?�������?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�������?�������?              �?      �?        333333�?�������?�$I�$I�?�m۶m��?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?I�$I�$�?۶m۶m�?      �?                      �?�j�j�j�?[�Z�Z��?�}ylE��?W'u_�?L�Ϻ��?�Y7�"��?      �?      �?]t�E�?t�E]t�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?                      �?��.���?t�E]t�?��8��8�?�q�q�?      �?      �?      �?        �������?�������?              �?      �?              �?              �?      �?              �?      �?        |���?>����?�������?ZZZZZZ�?�?�������?�$I�$I�?�m۶m��?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?      �?      �?      �?                      �?��}kdu�?�!H��h�?�{a���?a����?�q�q�?�q�q�?              �?�������?ZZZZZZ�?�a�a�?=��<���?      �?      �?              �?      �?        (�����?�5��P�?      �?      �?              �?      �?                      �?;�;��?vb'vb'�?�������?�������?�������?�������?      �?                      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�h
���?�_��e��?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJKc�HhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@>         ~                    �?�5�C��?H           ��@              A                    �?H��FG��?>           P~@               "       
             �?uvI��?�            �h@                                  �?�ȼB���?M            �[@                                 �]@�������?*             N@        ������������������������       �                     &@                      	          ����?����X�?"            �H@        ������������������������       �                     0@        	                           `@4���C�?            �@@        
                          �`@���Q��?             $@                     	          ����?؇���X�?             @       ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                  �a@�LQ�1	�?             7@                     
             �?��S���?
             .@        ������������������������       �                     @                                  �a@���!pc�?             &@                                   _@�q�q�?             @        ������������������������       �                     �?                                  g@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   @I@      �?              @                                   �F@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                !                   �x@`'�J�?#            �I@       ������������������������       �        "            �H@        ������������������������       �                      @        #       :                   �_@�H�a��?<            @U@        $       7       	          ����?�q���?             H@       %       2                    �?���|���?            �@@       &       /                    ]@�q�q�?             >@       '       (                   �Y@��.k���?	             1@        ������������������������       �                     @        )       .                    @K@և���X�?             ,@       *       -                    n@      �?             (@       +       ,                   �Z@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        0       1                   pc@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        3       6                    �?�q�q�?             @       4       5                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        8       9                    �?�r����?
             .@        ������������������������       �                      @        ������������������������       �        	             *@        ;       @       	             �?@-�_ .�?            �B@       <       =                   �b@������?             B@       ������������������������       �                    �@@        >       ?                   0c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        B       g       
             �?SSx~�?�            r@       C       X                    �?�Db�Aɵ?�            �n@       D       G                   �Z@�O���h�?o            �f@        E       F                   �Y@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        H       O                   Xp@`���i��?k             f@       I       N                    @J@����}��?J            �_@        J       M                    �?      �?             @@        K       L       	             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �        5            �W@        P       Q                    @M@��<D�m�?!            �H@       ������������������������       �                     A@        R       W                   �a@z�G�z�?             .@        S       V                    �O@���Q��?             @       T       U                   �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        Y       d                   �e@�U�=���?)            �P@       Z       c       	          ����?(;L]n�?&             N@        [       \                    �?�KM�]�?             3@        ������������������������       �                     �?        ]       b                    �L@�X�<ݺ?
             2@        ^       a                   @\@�����H�?             "@        _       `                    @K@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                    �D@        e       f                   �^@      �?             @       ������������������������       �                     @        ������������������������       �                     @        h       {                   Pd@��i#[�?             E@       i       x                    �?�d�����?             C@       j       u                   a@����X�?             <@       k       n       	             �?j���� �?
             1@        l       m                     P@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        o       p       	             �?z�G�z�?             $@        ������������������������       �                     @        q       r                    a@�q�q�?             @        ������������������������       �                     �?        s       t                    @N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        v       w                    d@�C��2(�?	             &@       ������������������������       �                     $@        ������������������������       �                     �?        y       z                    �G@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        |       }       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?               �       
             �?�?2����?
           {@        �       �                    �?���=��?g            @f@        �       �                   �c@�!���?             A@       �       �       	             �?j���� �?             1@       �       �                    �?r�q��?             (@       �       �                   �`@�C��2(�?             &@        �       �                   0l@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�IєX�?	             1@        �       �       	          `ff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        �       �                    �?ޚ)�?R             b@        �       �                    @J@r�qG�?             H@        ������������������������       �                     *@        �       �                    c@��
P��?            �A@        �       �       	          ����?"pc�
�?             &@       ������������������������       �                     @        �       �       	          hff@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    e@�q�q�?             8@       �       �                   `f@���!pc�?             6@       �       �                   �q@���N8�?             5@       �       �                    @�S����?             3@       �       �       
             �?և���X�?             @        ������������������������       �                      @        �       �       	          ����?���Q��?             @       �       �                   p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   P`@�q�Q�?9             X@        �       �                   �_@��V#�?            �E@       �       �                   pf@z�G�z�?            �A@       �       �                    �I@      �?             @@       �       �                   @Y@������?
             .@        ������������������������       �                     @        �       �                    @F@�8��8��?	             (@        �       �       	             �?      �?             @        ������������������������       �                      @        �       �                   0l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             1@        ������������������������       �                     @        �       �       
             �?      �?              @        ������������������������       �                     @        �       �       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?0��_��?            �J@       �       �       	          033�?6YE�t�?            �@@       �       �                   �r@�����H�?             ;@       �       �                   �h@$�q-�?             :@        ������������������������       �                     @        �       �                   �`@�KM�]�?             3@        ������������������������       �                     �?        �       �                    �?�X�<ݺ?             2@       ������������������������       �                     ,@        �       �                    �M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �Q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             4@        �       �       	             @�j�}��?�            �o@       �       �                   @g@0�`��!�?�            �o@       �       �                   �s@�I�?�_�?�            �o@       �       �                    c@0�M�n�?�             n@       �       �                    @L@������?�             l@       �       �                    �?�o"Q9a�?r            �f@       ������������������������       �        G             ]@        �       �                   Pc@��ɉ�?+            @P@        ������������������������       �                     �?        �       �                    �?     ��?*             P@        ������������������������       �        
             ,@        �       �                   c@p���?              I@        �       �                    �G@ �q�q�?             8@        �       �                   �[@ףp=
�?             $@        �       �                    Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@        ������������������������       �                     :@        �       �                    �L@�ʈD��?            �E@        �       �                    �?      �?             @        �       �                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?�?�|�?            �B@       ������������������������       �                     @@        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�t����?             1@        �       �                   0c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        
             ,@        �       �                   u@���!pc�?	             &@       �       �                    `@      �?             @        ������������������������       �                      @        �       �                    d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  G��*��?ܿ��j��?��)��?:D����?
^N��)�?��X��?5'��Ps�?3���+c�?�������?�������?              �?�$I�$I�?�m۶m��?              �?'�l��&�?m��&�l�?333333�?�������?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?d!Y�B�?Nozӛ��?�?�������?              �?F]t�E�?t�E]t�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?      �?      �?      �?                      �?      �?                      �?�?�������?              �?      �?        �������?TTTTTT�?�������?�������?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?�?�������?              �?�$I�$I�?۶m۶m�?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?        �؉�؉�?;�;��?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�?�������?      �?                      �?S�n0E�?к����?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?$�ɜoB�?�f�W�?�la�6ͦ?3��,��?������?�0&q��?�������?333333�?              �?      �?        F]t�E�?F]t�E�?�@ �?����~��?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?և���X�?��S�r
�?              �?�������?�������?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?e�M6�d�?�M6�d��?�?�������?(�����?�k(���?      �?        �q�q�?��8��8�?�q�q�?�q�q�?UUUUUU�?�������?              �?      �?                      �?              �?              �?      �?      �?              �?      �?        �<��<��?�a�a�?y�5���?Cy�5��?�$I�$I�?�m۶m��?ZZZZZZ�?�������?�m۶m��?�$I�$I�?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?F]t�E�?]t�E�?              �?      �?        �������?�������?      �?                      �?      �?      �?      �?                      �?���r�4�?��Ö�?���G?�?.p�\��?�������?�������?ZZZZZZ�?�������?UUUUUU�?�������?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?      �?              �?        �?�?UUUUUU�?UUUUUU�?              �?      �?              �?        ��8��8�?9��8���?�������?�������?      �?        PuPu�?_�_��?F]t�E�?/�袋.�?              �?�������?333333�?      �?                      �?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?�a�a�?��y��y�?(������?^Cy�5�?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?              �?      �?              �?              �?                      �?              �?              �?UUUUUU�?�������?6eMYS��?eMYS֔�?�������?�������?      �?      �?�?wwwwww�?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?      �?      �?                      �?              �?              �?      �?              �?      �?      �?              �?      �?              �?      �?        �V�9�&�?"5�x+��?e�M6�d�?'�l��&�?�q�q�?�q�q�?;�;��?�؉�؉�?              �?(�����?�k(���?      �?        �q�q�?��8��8�?              �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?              �?>>>>>>�?�?.Wr{�?'���H�?�i��i��?�eY�eY�?�����?�����?I�$I�$�?۶m۶m�?6��{��?�rS�<��?      �?        ?�?��? �����?              �?     ��?      �?      �?        \���(\�?{�G�z�?�������?UUUUUU�?�������?�������?      �?      �?      �?                      �?      �?              �?              �?        A_���?�}A_з?      �?      �?      �?      �?              �?      �?              �?        *�Y7�"�?к����?      �?        �������?�������?      �?                      �?<<<<<<�?�?UUUUUU�?UUUUUU�?      �?                      �?      �?        F]t�E�?t�E]t�?      �?      �?      �?              �?      �?              �?      �?              �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�:ohG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�=         �                    �?n�A��?H           ��@              =                    �?�<jV�?=           �~@               2                    �?�M�E$g�?{            �g@              1                    �?n�.P���?T             _@                                  �?P7Z�U��?J            �[@                                   b@���B���?             :@                                  �?���7�?             6@        ������������������������       �                     "@        	                           �D@$�q-�?	             *@        
                           _@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @               *                    �M@j���� �?8            @U@                                 �_@�ʻ����?.             Q@                                  f@��i#[�?             E@                                 h@��Sݭg�?            �C@        ������������������������       �                     ,@                                  �a@���Q��?             9@                     	             �?�θ�?	             *@                                 �^@r�q��?             (@                                  �L@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @               !                    U@$��m��?             :@                       
             �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        "       )       	             �?���!pc�?             6@       #       (       	          @33�?���N8�?             5@       $       %       
             �?�t����?             1@        ������������������������       �                     @        &       '                   �b@؇���X�?
             ,@       ������������������������       �        	             (@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        +       ,                   �h@�t����?
             1@        ������������������������       �                     @        -       .                    `P@؇���X�?             ,@       ������������������������       �                     &@        /       0                    �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             *@        3       <                    @M@      �?'             P@       4       7       
             �?��-�=��?            �C@        5       6                    ]@      �?             @       ������������������������       �                      @        ������������������������       �                      @        8       9                   Pj@ >�֕�?            �A@       ������������������������       �                     ?@        :       ;                     K@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     9@        >       U                    �?�/5mvq�?�             s@        ?       B                    @I@�^�����?            �E@        @       A       	              @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        C       P                   hu@���@��?            �B@       D       O                    �?6YE�t�?            �@@       E       H                   `^@�q�q�?             8@        F       G                   `c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        I       L       	          033�?R���Q�?             4@       J       K       
             �?�IєX�?	             1@       ������������������������       �                     0@        ������������������������       �                     �?        M       N                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        Q       T       
             �?      �?             @       R       S                   �w@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        V       y       
             �? 	��p�?�            Pp@       W       t                    �? \sF��?�            @l@       X       s                    �?��Ͻ��?n            @e@       Y       Z                   �U@`�BX�l�?W             a@        ������������������������       �                     �?        [       \       
             �?�IєX�?V             a@        ������������������������       �        
             1@        ]       b                    �?T(y2��?L            �]@        ^       a                     G@ 7���B�?             ;@        _       `       	             @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     9@        c       d                   e@�c:��?:             W@        ������������������������       �                     :@        e       r                   0c@��IF�E�?+            �P@       f       q       	          ����?     p�?*             P@        g       j                   0i@$G$n��?            �B@        h       i                    �C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        k       p                   �Z@�g�y��?             ?@        l       o                   `a@؇���X�?             @        m       n                    Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                     ;@        ������������������������       �                      @        ������������������������       �                    �@@        u       x                   �i@�h����?#             L@        v       w                   `X@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                    �C@        z       �                    �?4�2%ޑ�?            �A@       {       |                   ``@��+7��?             7@        ������������������������       �                     $@        }       ~                   �h@��
ц��?
             *@        ������������������������       �                     @               �                    �L@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �       	             �?r�q��?             (@       ������������������������       �                     @        �       �       	             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	             �?����'�?           �z@       �       �                    �?h8"J{�?�            �r@       �       �                    �? �\���?[            �c@        �       �                    �?��2(&�?             6@       �       �                    �?r�q��?             2@        ������������������������       �                     �?        �       �                   �a@�t����?
             1@       ������������������������       �                     .@        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?�?�0�!�?O             a@        �       �                    �?�eP*L��?             &@       �       �                   �_@���Q��?             $@        ������������������������       �                     @        �       �                     C@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        G            @_@        �       �                    �?d}h���?Z            �a@       �       �       
             �?r�q��?G             [@        �       �                   b@     ��?             @@        ������������������������       �                     *@        �       �                    @B@�d�����?             3@        ������������������������       �                     �?        �       �                   �l@�<ݚ�?             2@        ������������������������       �                     "@        �       �                   Pc@X�<ݚ�?             "@       �       �                   Pm@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        1             S@        �       �       
             �?      �?             @@        �       �                    �?z�G�z�?	             .@        �       �                    `P@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �        
             1@        �       �                    �?     ��?V             `@        �       �       
             �?�חF�P�?             ?@       �       �                    �?�E��ӭ�?             2@        ������������������������       �                     @        �       �                    @�eP*L��?	             &@       �       �       	          ����?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             *@        �       �                    @F@��Lz���??            @X@        �       �       	          033@���!pc�?             &@       �       �                    @B@�����H�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�a7���?7            �U@       �       �                    �M@����"�?"             M@       �       �                    �?����X�?             E@        �       �                    �K@��S���?             .@        ������������������������       �                     @        �       �                    @z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        �       �                    e@�+$�jP�?             ;@       �       �                   @Z@�LQ�1	�?             7@        �       �       	          ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �^@ףp=
�?             4@        �       �       	             �?�q�q�?             @       �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   Pi@�IєX�?             1@       �       �                   @c@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    U@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?      �?             0@        �       �       	          `ff�?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �j@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   pb@��X��?             <@       �       �       
             �?z�G�z�?             4@       �       �                   �X@�	j*D�?             *@        ������������������������       �                     �?        �       �       	          ���@      �?             (@       �       �                   �`@�����H�?	             "@        �       �                    ]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �K@�q�q�?             @        ������������������������       �                     �?        �       �       	          `ff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                     P@      �?              @       �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  >��=���?a�a��?鰑�?<�œ[<�?���Q���?� &W��?�9�s��?c�1�c�?Nq��$�?c��2��?��؉���?ى�؉��?�.�袋�?F]t�E�?      �?        �؉�؉�?;�;��?      �?      �?              �?      �?              �?                      �?ZZZZZZ�?�������?<<<<<<�?�������?�<��<��?�a�a�?�i�i�?�|˷|��?              �?�������?333333�?ى�؉��?�؉�؉�?�������?UUUUUU�?]t�E�?F]t�E�?      �?                      �?              �?              �?              �?      �?        �N��N��?vb'vb'�?      �?      �?              �?      �?        F]t�E�?t�E]t�?�a�a�?��y��y�?�������?�������?              �?۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?�������?�������?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?�A�A�?}˷|˷�?      �?      �?              �?      �?        �A�A�?��+��+�?              �?      �?      �?      �?                      �?              �?������?�k(����?֔5eMY�?�5eMYS�?�������?UUUUUU�?      �?                      �?к����?L�Ϻ��?e�M6�d�?'�l��&�?�������?UUUUUU�?      �?      �?      �?                      �?333333�?333333�?�?�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �{a���?������?Vzja���?[X驅��?�?NNNNNN�?��;�HѰ?�������?      �?        �?�?              �?�5�5�?�F��F��?h/�����?	�%����?      �?      �?              �?      �?                      �?8��Moz�?Y�B���?              �?'�l��&�?�l��&��?      �?     ��?���L�?к����?UUUUUU�?UUUUUU�?              �?      �?        �B!��?��{���?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?              �?              �?      �?                      �?�$I�$I�?۶m۶m�?�?�?      �?                      �?              �?�A�A�?�������?Y�B��?zӛ����?              �?�؉�؉�?�;�;�?              �?      �?      �?      �?                      �?UUUUUU�?�������?              �?�������?333333�?      �?                      �?�b���i�?�u&`�X�?Y���a��?���DxR�?���7a�?�3���?��.���?t�E]t�?�������?UUUUUU�?              �?<<<<<<�?�?      �?                      �?      �?        �������?�����Ң?t�E]t�?]t�E�?333333�?�������?              �?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?        I�$I�$�?۶m۶m�?�������?UUUUUU�?      �?      �?              �?Cy�5��?y�5���?              �?9��8���?�q�q�?      �?        r�q��?�q�q�?�������?UUUUUU�?              �?      �?                      �?      �?              �?      �?�������?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?             @�?     ��?�Zk����?��RJ)��?�q�q�?r�q��?      �?        t�E]t�?]t�E�?      �?      �?              �?      �?              �?              �?        Z�D�a��?Ӱ�,O"�?F]t�E�?t�E]t�?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�qG��?qG�w�?�i��F�?	�=����?�$I�$I�?�m۶m��?�������?�?      �?        �������?�������?              �?      �?        B{	�%��?/�����?Y�B��?��Moz��?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?�?�?      �?      �?              �?      �?                      �?      �?      �?              �?      �?              �?      �?      �?      �?      �?                      �?      �?      �?      �?                      �?%I�$I��?n۶m۶�?�������?�������?;�;��?vb'vb'�?      �?              �?      �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�RrhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK녔h��B�:         �       	          033�?V�2���?A           ��@              a                    �?>��"��?B           8�@                                 �O@��ʙ�5�?           0z@                                   �?D>�Q�?%             J@                      	          ����?�û��|�?             7@                                 �Y@@�0�!��?             1@        ������������������������       �                     �?               	                    �?      �?             0@       ������������������������       �                      @        
              	          �����      �?              @        ������������������������       �                     �?                                  0a@؇���X�?             @                                   \@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     =@                                    �?�������?�            �v@                                  Pt@�h����?D             \@                                  `@@䯦s#�??            �Z@       ������������������������       �        %             P@                                   �?�Ń��̧?             E@                                   �K@ףp=
�?             $@       ������������������������       �                      @                                  �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@                                   �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        !       2       
             �?������?�            �o@        "       1                   0f@@�r-��?            �M@       #       &                    �E@���5��?            �L@        $       %                   �_@      �?              @       ������������������������       �                     @        ������������������������       �                     @        '       .                    @��<D�m�?            �H@       (       )       	          ����?`�q�0ܴ?            �G@       ������������������������       �                     E@        *       -                    �?���Q��?             @       +       ,                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        /       0                     O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        3       \                    �O@�)���Y�?}            �h@       4       S                   �b@ ��@��?x            `g@       5       B                    �?�1��?o            �e@        6       7                    �E@�t����?             A@        ������������������������       �                     (@        8       9                   �e@"pc�
�?             6@        ������������������������       �                     �?        :       A                    �?؇���X�?             5@        ;       @                   �d@և���X�?             @       <       ?       	          ����?      �?             @       =       >                   pn@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             ,@        C       H                    Z@�|y���?Z            `a@        D       E                    �J@      �?              @       ������������������������       �                     @        F       G                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        I       P       	          833�?@��A1ʞ?U            ``@       J       O                   pi@ >��@�?R            @_@        K       L                    @N@�Ń��̧?             E@       ������������������������       �                     C@        M       N                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        :            �T@        Q       R                     @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        T       Y                    �J@և���X�?	             ,@       U       X                    �D@      �?              @        V       W                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Z       [                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ]       `                   �a@X�<ݚ�?             "@       ^       _                   �j@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        b       s       
             �?��:M�?>             Y@       c       r                   `f@lGts��?#            �K@       d       e                    l@h�WH��?"             K@       ������������������������       �                     <@        f       o                    �O@���B���?             :@       g       h                    \@؇���X�?             5@        ������������������������       �                     �?        i       l                    �F@ףp=
�?             4@        j       k       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        m       n                   �l@�X�<ݺ?
             2@        ������������������������       �                     �?        ������������������������       �        	             1@        p       q                    @P@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        t       �                   Pd@���Q��?            �F@       u       v                    �?�eP*L��?            �@@        ������������������������       �                     @        w       �                    �?���Q��?             >@       x                           I@$��m��?             :@        y       ~       	             �?r�q��?             (@       z       {                   �a@����X�?             @        ������������������������       �                     @        |       }                    [@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �c@      �?
             ,@       �       �                    �K@�<ݚ�?             "@       ������������������������       �                     @        �       �                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?V�s	J��?�            �x@        �       �                   Xr@b��虠�?W            `a@       �       �                    �?�������?H            @\@        �       �       
             �?�d�����?             3@        ������������������������       �                     @        �       �                   �Z@��S�ۿ?             .@        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   0`@�*/�8V�?:            �W@        �       �                    �Q@ 	��p�?             =@       ������������������������       �                     :@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�4��?(            @P@       �       �                    �?��+��?            �B@        �       �                   pb@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          ���
@*;L]n�?             >@       �       �       	             @      �?             :@       �       �       
             �?�����?             3@       �       �                   �\@�eP*L��?             &@        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                     @        �       �       	          `ff�?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?؇���X�?             <@        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �L@�8��8��?             8@        �       �                    �K@"pc�
�?             &@       �       �                    �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     *@        �       �                    �?$�q-�?             :@        ������������������������       �                     *@        �       �                     L@8�Z$���?             *@       ������������������������       �                     $@        �       �       
             �?�q�q�?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �e@$�q-�?�            @p@        �       �                    @M@�(\����?0             T@        ������������������������       �                     B@        �       �                   P`@���7�?             F@       ������������������������       �                    �C@        �       �                    �?���Q��?             @       �       �                    �?      �?             @       �       �       	             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?ףp=
�?x            �f@       �       �                   �f@˒�#�?g            �b@        ������������������������       �                     �?        �       �                   Pj@@9G��?f            `b@        �       �                   �\@�LQ�1	�?             7@        ������������������������       �                     @        ������������������������       �                     4@        �       �                     R@�â��,�?V             _@       �       �                    `@p�,�V��?T            @^@        ������������������������       �                     D@        �       �                    �?F|/ߨ�?;            @T@        �       �                   ``@؇���X�?             ,@        ������������������������       �                     �?        �       �                   p`@$�q-�?             *@        �       �                   �^@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �        /            �P@        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?     ��?             @@       �       �                    `P@�G��l��?             5@       �       �       	          ����?ҳ�wY;�?
             1@       �       �                   �q@d}h���?             ,@       ������������������������       �                     $@        �       �                   �r@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  � ���Y�?�o�6S�?�����?��R�O2�?9����^�?����B�?vb'vb'�?b'vb'v�?��,d!�?8��Moz�?�������?ZZZZZZ�?      �?              �?      �?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?�ɑA~��?�ٸ�j�?۶m۶m�?�$I�$I�?R����?�x+�R�?      �?        ��<��<�?�a�a�?�������?�������?      �?              �?      �?      �?                      �?      �?        �������?UUUUUU�?              �?      �?        wwwwww�?�?��c+���?'u_�?��Gp�?�}��?      �?      �?              �?      �?        և���X�?��S�r
�?W�+�ɥ?��F}g��?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?              �?        Dc}h��?������?��:����?�)��˱?��#���?+���}��?<<<<<<�?�?      �?        /�袋.�?F]t�E�?              �?۶m۶m�?�$I�$I�?�$I�$I�?۶m۶m�?      �?      �?      �?      �?      �?                      �?              �?      �?              �?        ���1O�?'!����?      �?      �?      �?              �?      �?              �?      �?        �ֆi��?qBJ�eD�?X9��v��?����Mb�?��<��<�?�a�a�?      �?              �?      �?      �?                      �?      �?        �������?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?              �?      �?        �q�q�?r�q��?UUUUUU�?�������?      �?                      �?      �?        ��Q��?q=
ףp�?�־a�?�<%�S��?B{	�%��?��^B{	�?              �?ى�؉��?��؉���?�$I�$I�?۶m۶m�?      �?        �������?�������?      �?      �?              �?      �?        �q�q�?��8��8�?      �?                      �?�������?333333�?      �?                      �?      �?        333333�?�������?]t�E�?t�E]t�?      �?        �������?333333�?vb'vb'�?�N��N��?UUUUUU�?�������?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?              �?        䤑�FN�?ǖ[nl�?�j����?������?�ZX驅�?��S+=�?Cy�5��?y�5���?              �?�������?�?              �?      �?        AL� &W�?�٨�l��?�{a���?������?              �?UUUUUU�?UUUUUU�?              �?      �?        �Z��Z��?�R+�R+�?*�Y7�"�?�S�n�?�$I�$I�?۶m۶m�?              �?      �?        """"""�?�������?      �?      �?Q^Cy��?^Cy�5�?]t�E�?t�E]t�?              �?�m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?F]t�E�?/�袋.�?�������?�������?      �?                      �?      �?                      �?�؉�؉�?;�;��?      �?        ;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?;�;��?�؉�؉�?�������?333333�?              �?F]t�E�?�.�袋�?              �?�������?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?        �������?�������?v�)�Y7�?�g�`�|�?      �?        9/���?������?Y�B��?��Moz��?      �?                      �?�c�1Ƙ?:�s�9�?���k��?ˠT�x�?              �?�����H�?�Hx�5�?�$I�$I�?۶m۶m�?      �?        ;�;��?�؉�؉�?      �?      �?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?1�0��?��y��y�?�������?�������?I�$I�$�?۶m۶m�?      �?              �?      �?              �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJF�yhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKh��B�;         �       	          033�?���3L�?L           ��@              I                    �?Z�ݓ�?E           (�@                                   �?j$ޗQ�?�            �i@                                   �M@�z�G��?             >@                                  �?�q�q�?             8@                                 �T@��2(&�?             6@        ������������������������       �                     �?               	                    �?�����?             5@       ������������������������       �        	             .@        
                           �?�q�q�?             @        ������������������������       �                      @                                  `r@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                                  �\@�q�q�?             @        ������������������������       �                     �?                                   e@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?               @                    �?H��Q6�?t            �e@                     
             �?U��K��?Q            @^@                                    M@@4և���?$             L@       ������������������������       �                     @@                                  �l@r�q��?             8@                                 �k@���N8�?             5@       ������������������������       �                     2@                                  �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                1                   pc@�7�֥��?-            @P@       !       .                    @O@R���Q�?             D@       "       #                    ]@������?            �B@        ������������������������       �                     @        $       +                   @E@�r����?             >@        %       (                    �?և���X�?             @        &       '       	             �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        )       *                    `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ,       -                    �?�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        /       0                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        2       ?                    �? �o_��?             9@       3       6                   �d@��S���?             .@        4       5                    �C@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        7       8                   Pe@�q�q�?             "@        ������������������������       �                     @        9       <                    �?      �?             @       :       ;                   f@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        =       >                    �D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        A       B                    k@0��_��?#            �J@       ������������������������       �                    �B@        C       D       
             �?     ��?             0@       ������������������������       �                     "@        E       H                   ``@����X�?             @        F       G                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        J       W                   `@H6���r�?�            �s@        K       L       
             �?R_u^|�?)            �Q@        ������������������������       �                    �B@        M       N                    �?l��\��?             A@        ������������������������       �                     &@        O       T                    q@�LQ�1	�?             7@       P       Q                    _@�}�+r��?             3@       ������������������������       �                     0@        R       S                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        U       V                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        X       q       
             �?�y)|���?�            @n@        Y       p                   xq@��6���?             E@       Z       [                   �Q@�xGZ���?            �A@        ������������������������       �                     @        \       e                   `m@���@M^�?             ?@        ]       d                   0m@8�Z$���?	             *@       ^       c                    �?�<ݚ�?             "@       _       `                   �c@      �?              @        ������������������������       �                     @        a       b                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        f       g                   �m@X�<ݚ�?	             2@        ������������������������       �                     @        h       o                    �?և���X�?             ,@       i       n                    �?�����H�?             "@       j       m       	          ����?؇���X�?             @        k       l                     E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        r       y                    �L@`2U0*��?{             i@       s       t                    �J@������?e            `d@       ������������������������       �        P             `@        u       x                    �?��?^�k�?            �A@        v       w                   �o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @@        z                          �s@��G���?            �B@       {       |       	          833�?ףp=
�?             >@       ������������������������       �                     8@        }       ~                     O@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �       	          ����?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�ij�?           y@        �       �                   �a@B�
k���?/            �P@       �       �       	          pff�?f.i��n�?!            �F@       �       �       
             �?     ��?             @@        ������������������������       �                     �?        �       �                   �_@��� ��?             ?@        ������������������������       �                     (@        �       �                    �?���y4F�?             3@       �       �                    �K@��S�ۿ?
             .@       ������������������������       �                     $@        �       �                    �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �                    �I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�	j*D�?             *@       ������������������������       �                     "@        ������������������������       �                     @        �       �                   �c@"pc�
�?             6@       �       �                    @H@�KM�]�?             3@        �       �                   Xs@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             ,@        �       �                   �d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@�>q���?�            �t@       �       �       	          ����?�~�H��?�            pp@        �       �                    �?��s����?%            �O@       �       �                   �[@���y4F�?             �L@        ������������������������       �                     &@        �       �                    �?��+7��?             G@        �       �                    @I@      �?             0@        ������������������������       �                     @        �       �                   `@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                    �K@��S�ۿ?             >@       ������������������������       �                     4@        �       �                   @_@z�G�z�?             $@       �       �                    �?�����H�?             "@        ������������������������       �                      @        �       �                   �]@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?DGr���?�             i@       �       �       	          ����?ܷ��?��?^             b@        �       �                    �?*
;&���?             G@       ������������������������       �                     ;@        �       �                   �l@p�ݯ��?	             3@       �       �       
             �?���|���?             &@       �       �                   �j@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �F@�"P��?C            �X@        �       �                    �?�q�q�?
             .@        ������������������������       �                     @        �       �                   �r@r�q��?             (@       �       �                   �i@�C��2(�?             &@       ������������������������       �                      @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �J@h�����?9             U@        �       �                    @J@ףp=
�?             4@       ������������������������       �                     .@        �       �                   @]@���Q��?             @       �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �       
             �?     ��?*             P@       ������������������������       �        %             K@        �       �                   �`@ףp=
�?             $@        �       �                   `^@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          pff@h㱪��?(            �K@       ������������������������       �                      G@        �       �                   �c@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                    c@$]��<C�?-            �Q@       �       �                    �?Xny��?'            �N@       �       �                    @Q@`Ӹ����?            �F@       ������������������������       �                    �E@        ������������������������       �                      @        �       �                    @I@     ��?
             0@        ������������������������       �                     @        �       �                    `P@      �?             $@       �       �                    �L@����X�?             @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �       	          hff@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �t�b�b6     h�h)h,K ��h.��R�(KK�KK��hb�B�  &���^B�?�%���^�?�J�_�?�uj��@�?FFFFFF�?�������?ffffff�?333333�?UUUUUU�?�������?��.���?t�E]t�?              �?=��<���?�a�a�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        �@&�d�?��l���?*L�9��?��!pc�?�$I�$I�?n۶m۶�?              �?UUUUUU�?�������?�a�a�?��y��y�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �B/�B/�?z�z��?333333�?333333�?��g�`��?к����?      �?        �������?�?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?�Mozӛ�?d!Y�B�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �Q����?
ףp=
�?�������?�?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�V�9�&�?"5�x+��?              �?      �?      �?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UX4���?«�.��?2~�ԓ��?�@�6�?              �?------�?�������?      �?        ��Moz��?Y�B��?�5��P�?(�����?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        &ޏ���?�g���e�?=��<���?b�a��?�_�_�?�A�A�?              �?�s�9��?�c�1��?;�;��?;�;��?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �q�q�?r�q��?              �?�$I�$I�?۶m۶m�?�q�q�?�q�q�?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?                      �?              �?���Q��?{�G�z�?<^l	���?)��I� y?      �?        _�_��?�A�A�?UUUUUU�?UUUUUU�?      �?                      �?      �?        #�u�)��?v�)�Y7�?�������?�������?      �?              �?      �?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        |��O���?��,���?L�*g��?g��1��?�`�`�?�>�>��?      �?      �?              �?�{����?�B!��?      �?        6��P^C�?(������?�������?�?      �?        �������?�������?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?;�;��?vb'vb'�?              �?      �?        F]t�E�?/�袋.�?(�����?�k(���?�������?333333�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?qZ�}�z�?d)�`W��?���-g:�?�H�x�?�a�a�?z��y���?(������?6��P^C�?              �?Y�B��?zӛ����?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �?�������?              �?�������?�������?�q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?              �?      �?              �?                      �?��(\�µ?H�z�G�?a���{�?��=���?8��Moz�?���,d!�?              �?Cy�5��?^Cy�5�?]t�E]�?F]t�E�?333333�?�������?              �?      �?              �?                      �?[�R�֯�?��+j�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?�������?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �$I�$I�?�m۶m��?�������?�������?              �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?     ��?              �?�������?�������?      �?      �?              �?      �?                      �?��)A��?־a���?              �?�q�q�?9��8���?              �?      �?        �'�K=�?6���?�}�K�`�?C��6�S�?l�l��??�>��?              �?      �?              �?      �?              �?      �?      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?ffffff�?333333�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJܓ�!hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KKh��B�;         �                    �?��+�?E           ��@              !                    �?�ns��#�?=           P@                                  �a@�\����?+            �P@                                  �?���|���?             F@                     
             �?p9W��S�?             C@                                  �?j���� �?             1@                                  �p@      �?              @       ������������������������       �                     @        	       
                   �t@      �?             @        ������������������������       �                     @        ������������������������       �                     �?                                  �g@�<ݚ�?             "@        ������������������������       �                     �?                                   �O@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                   �?���N8�?             5@                                   `@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             2@                                  �[@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                      	          ����?�X����?             6@                                  Pd@      �?              @        ������������������������       �                      @        ������������������������       �                     @                                    �H@@4և���?             ,@                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             (@        "       I                    @H@P��ʹ�?           0{@        #       8       
             �?�n����?@            @Z@       $       %                    @D@ >�֕�?)            �Q@        ������������������������       �                     :@        &       -                    �?�C��2(�?             F@        '       ,                    �?�r����?	             .@       (       +                    �E@"pc�
�?             &@        )       *                    \@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        .       5                   pb@ 	��p�?             =@       /       0       	             �? 7���B�?             ;@       ������������������������       �        	             2@        1       4                   �h@�����H�?             "@        2       3                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        6       7                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        9       H                    �?<=�,S��?            �A@       :       =                    �?¦	^_�?             ?@        ;       <                    @F@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        >       E                   �b@r�q��?             8@       ?       B                    �?ףp=
�?             4@       @       A                   �_@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@        C       D                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        F       G                   po@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        J       e       
             �?t���|�?�            �t@       K       b                   pz@`2U0*��?�            @o@       L       a                    �?��d�?�             o@       M       \                    �O@p��D׀�?j            �c@       N       [                   �m@���U�?Q            �\@       O       X                   �c@�FVQ&�?4            �P@       P       W                    �K@�i�y�?2            �O@        Q       T                   Pl@�>����?             ;@       R       S                   �W@ �q�q�?             8@        ������������������������       �                     �?        ������������������������       �                     7@        U       V                     J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     B@        Y       Z                   �d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     H@        ]       `       	          `ff�?�Ra����?             F@        ^       _                   �[@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                    �@@        ������������������������       �        8            �V@        c       d       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       {                    �?��Q���?.             T@        g       v                    �?��+��?            �B@       h       o       	            �?�f7�z�?             =@       i       n                    b@���y4F�?             3@       j       m                   �q@r�q��?
             2@       k       l                    V@      �?	             0@        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                      @        ������������������������       �                     �?        p       u                   �s@z�G�z�?             $@       q       t                   `a@�����H�?             "@        r       s                   @a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        w       x                   ``@      �?              @       ������������������������       �                     @        y       z                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        |       �                    p@RB)��.�?            �E@       }       �                   �^@<���D�?            �@@        ~              	             �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                     M@ 7���B�?             ;@        �       �                    @L@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             6@        �       �                   �r@      �?             $@        �       �       	          ����?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?&���v�?           z@        �       �                   �c@     ��?c             d@       �       �                   p`@<�I<���?N             `@       �       �                   P`@h��@D��?)            �Q@        �       �                   �s@@�0�!��?             A@       �       �                     N@6YE�t�?            �@@       �       �                    �?�GN�z�?             6@       �       �                    �K@�t����?             1@       �       �                   �_@؇���X�?             ,@       ������������������������       �                     "@        �       �                    �J@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �?�?�|�?            �B@        �       �                   c@�����H�?             "@       ������������������������       �                     @        �       �                   @e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     <@        �       �                    @E@8^s]e�?%             M@        ������������������������       �                     @        �       �                   o@������?#             K@       �       �                   Pk@���@M^�?             ?@       �       �                   �a@      �?             0@        �       �                   �W@z�G�z�?             @        �       �                    a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �       	          `ff@������?
             .@       �       �                    �?8�Z$���?	             *@        ������������������������       �                     �?        �       �                   �m@�8��8��?             (@       ������������������������       �                     @        �       �                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �e@���}<S�?             7@       �       �                   �b@�}�+r��?             3@       ������������������������       �                     (@        �       �                   0c@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?f���M�?             ?@        �       �                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                   p@      �?             4@       �       �                   pm@����X�?
             ,@       �       �                    �?      �?              @        ������������������������       �                     @        �       �                   �[@z�G�z�?             @        �       �                   �d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �]@�"��#�?�            p@        �       �                   `\@      �?             D@       ������������������������       �                     @@        �       �       	             �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   `Q@����Ձ�?�             k@        �       �                   `_@�z�G��?             $@        ������������������������       �                      @        �       �                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�n����?�            �i@       �       �                    @L@�?�|�?v             g@       ������������������������       �        `             c@        �       �                    �M@6YE�t�?            �@@        �       �       	          @33�?�q�q�?             (@       �       �                    �?�<ݚ�?             "@       �       �                    @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        �       �                    �?�C��2(�?             6@        �       �       	             �?�q�q�?             @       �       �                   Pd@���Q��?             @       �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  f�,I��?Ͱ�w[��?�C�e�	�?/�����?���>��?>����?]t�E]�?F]t�E�?�k(����?l(�����?ZZZZZZ�?�������?      �?      �?      �?              �?      �?              �?      �?        �q�q�?9��8���?      �?              �?      �?              �?      �?        ��y��y�?�a�a�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?      �?                      �?]t�E]�?�E]t��?      �?      �?              �?      �?        �$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?^�(ٵ��?)ٵ��]�? �����?8�8��?�A�A�?��+��+�?              �?F]t�E�?]t�E�?�?�������?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�{a���?������?h/�����?	�%����?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?�A�A�?X|�W|��?��Zk���?�RJ)���?�$I�$I�?�m۶m��?              �?      �?        �������?UUUUUU�?�������?�������?�?�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?              �?      �?                      �?��?����?j�ƀi�?{�G�z�?���Q��?�RJ)���?�Zk����?T:�g *�?[܄�]-�?p�}��?	�#����?|���?>����?AA�?�������?h/�����?�Kh/��?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?]t�E�?]t�E]�?]t�E�?t�E]t�?              �?      �?                      �?              �?      �?      �?      �?                      �?�������?333333�?*�Y7�"�?�S�n�?O#,�4��?a���{�?6��P^C�?(������?�������?UUUUUU�?      �?      �?              �?      �?                      �?              �?�������?�������?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?              �?      �?              �?      �?      �?      �?                      �?���)k��?S֔5eM�?|���?|���?      �?      �?              �?      �?        h/�����?	�%����?�������?�������?              �?      �?                      �?      �?      �?�������?UUUUUU�?      �?                      �?              �?_�Q�#�?C�\ɸ��?      �?      �?4�9c��?sƜ1g��?�'�K=�?��V��?�������?ZZZZZZ�?e�M6�d�?'�l��&�?]t�E�?�袋.��?�������?�������?�$I�$I�?۶m۶m�?              �?�������?333333�?      �?                      �?      �?                      �?              �?      �?        к����?*�Y7�"�?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?	�=����?|a���?      �?        {	�%���?B{	�%��?�c�1��?�s�9��?      �?      �?�������?�������?      �?      �?              �?      �?                      �?              �?wwwwww�?�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?                      �?              �?d!Y�B�?ӛ���7�?(�����?�5��P�?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?      �?      �?                      �?��RJ)��?��Zk���?]t�E�?F]t�E�?      �?                      �?      �?      �?�m۶m��?�$I�$I�?      �?      �?      �?        �������?�������?      �?      �?      �?                      �?              �?      �?                      �?�!�!�!�?���?      �?      �?      �?              �?      �?      �?                      �?��}��?�`^0/��?ffffff�?333333�?              �?      �?      �?      �?                      �?�<����?j6��bP�?*�Y7�"�?к����?      �?        '�l��&�?e�M6�d�?�������?�������?9��8���?�q�q�?�m۶m��?�$I�$I�?      �?                      �?      �?                      �?      �?        ]t�E�?F]t�E�?UUUUUU�?UUUUUU�?333333�?�������?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��]hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@=         �                    �?�O(�.��?E           ��@              s                    �?�qi�-}�?C           �@              4                    �?ܚ�R��?�             w@               +                    �?�Z����?V             a@                     
             �?��J�fj�?G            �[@                                 �]@&y�X���?&             M@        ������������������������       �        
             0@                                   b@0,Tg��?             E@        	                          �u@�q�q�?             8@       
                           �?      �?             4@        ������������������������       �                     "@                                  0`@�C��2(�?             &@        ������������������������       �                     @                                   p@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                  `]@�X�<ݺ?             2@                      	          @33�?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             &@               *       	          ����?�q����?!            �J@              !                    �?`�Q��?             I@                                   d@������?
             1@                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     @                                    �I@�C��2(�?             &@                                   \@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        "       )                   �^@�C��2(�?            �@@       #       (                   @^@@�0�!��?             1@       $       %                   pl@��S�ۿ?
             .@       ������������������������       �                      @        &       '                   �b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             0@        ������������������������       �                     @        ,       3       	             �?ȵHPS!�?             :@       -       2                    T@ �q�q�?             8@        .       /       
             �?      �?             @        ������������������������       �                     �?        0       1                     H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        
             4@        ������������������������       �                      @        5       h                   pb@\�#���?�            �l@       6       _       	          ����?`�H�/��?�            �i@       7       L                    �?�X�C�?G             \@       8       E                   �_@�gc� �?4            �T@       9       D       	          ����?@4և���?#             L@        :       C                    �O@"pc�
�?             6@       ;       @       
             �?؇���X�?             5@       <       ?                   @\@�X�<ݺ?
             2@        =       >       	             �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        A       B                     M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        F       I                   pb@�<ݚ�?             ;@       G       H       	          ����?�}�+r��?             3@       ������������������������       �        
             2@        ������������������������       �                     �?        J       K                    @J@      �?              @        ������������������������       �                     @        ������������������������       �                     @        M       X                   ``@�c�Α�?             =@       N       O                   �W@և���X�?
             ,@        ������������������������       �                      @        P       W                     O@      �?	             (@       Q       T                    @L@���Q��?             $@        R       S                    ^@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        U       V                   �Y@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Y       ^                   �s@�r����?	             .@       Z       ]                   @U@@4և���?             ,@        [       \       	             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        `       a                    �?��<b�ƥ?@             W@        ������������������������       �                      @        b       c                   �W@����?�?>            �V@        ������������������������       �                     �?        d       e                   �`@ }�Я��?=            @V@       ������������������������       �        +             P@        f       g                    U@`2U0*��?             9@        ������������������������       �                     �?        ������������������������       �                     8@        i       l                   pn@�5��?             ;@        j       k                   �i@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        m       r                    �?      �?	             0@        n       q       	          `ff�?����X�?             @       o       p                   �e@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        t       w                   �Q@�nkK�?W            @a@        u       v                   Pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        x       y       	          ����?�?�0�!�?U             a@        ������������������������       �                     B@        z       �                    �R@P���Q�??             Y@       {       �       	          833�?`�(c�?>            �X@        |       }                    �G@�z�G��?             $@        ������������������������       �                     @        ~                          �b@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        7             V@        ������������������������       �                      @        �       �                    �?��m�_�?           �y@       �       �                   `Q@��֩�X�?�            �u@        �       �                    �?�n_Y�K�?             :@       �       �       
             �?�d�����?             3@       �       �                    `Q@��S�ۿ?
             .@       ������������������������       �        	             ,@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          `ff�?\���(\�?�             t@       �       �                   �l@��a��?�            @n@        �       �                   �]@ ��7��?G            �^@        �       �                    �?�nkK�?             7@       ������������������������       �                     1@        �       �                   �d@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        8            �X@        �       �                   �g@2Tv���?L             ^@       �       �                    @|�9ǣ�?K            �]@       �       �                   @m@�>����?E             [@        �       �                   pe@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?`'�J�?B            �Y@       �       �       
             �?@�E�x�??            �X@        �       �                    @L@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �G@�|���?9             V@        �       �                     G@P�Lt�<�?             C@       ������������������������       �                     B@        �       �                    o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     I@        �       �                   �c@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    b@�z�G��?             $@       �       �                   �p@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �       	          033�?�n_Y�K�?/            �S@       �       �                    �L@�k��(A�?"            �M@       �       �                   �f@R���Q�?             D@        ������������������������       �                      @        �       �                   �l@�KM�]�?             C@        ������������������������       �        	             2@        �       �                    �?z�G�z�?             4@       �       �                   @_@@4և���?             ,@        �       �       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                   �l@      �?             @        ������������������������       �                     �?        �       �                    @L@���Q��?             @       �       �       
             �?      �?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@D�n�3�?
             3@       �       �       	          `ff�?և���X�?             ,@       �       �                    �R@�q�q�?             "@       �       �                     N@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�����?             3@        ������������������������       �                     @        �       �       
             �?     ��?
             0@        ������������������������       �                      @        �       �                   ``@@4և���?	             ,@        �       �                   @_@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?-            �P@       �       �                    �?�^�����?            �E@        ������������������������       �                      @        �       �                   �X@<=�,S��?            �A@        ������������������������       �                     �?        �       �                   �`@ҳ�wY;�?             A@        �       �                   �k@"pc�
�?             &@       ������������������������       �                      @        �       �                    [@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@�LQ�1	�?             7@        ������������������������       �                     @        �       �       
             �?r�q��?             2@        �       �                   �d@      �?             @        ������������������������       �                      @        �       �                   �^@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             (@        �       �       	          @33�?�LQ�1	�?             7@        �       �       
             �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �\@�X�<ݺ?             2@        �       �       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             .@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �6S���?��rV��?����Q�?MĖ��+�?����7��?���,d!�?��s2}��?�J���?к����?�"�u�)�?�i��F�?��FX��?              �?1�0��?�y��y��?�������?�������?      �?      �?      �?        F]t�E�?]t�E�?              �?�������?�������?              �?      �?                      �?�q�q�?��8��8�?�$I�$I�?۶m۶m�?              �?      �?                      �?�Cj��V�?�x+�R�?��(\���?{�G�z�?�?xxxxxx�?      �?      �?      �?                      �?F]t�E�?]t�E�?�������?�������?              �?      �?                      �?]t�E�?F]t�E�?ZZZZZZ�?�������?�������?�?      �?        ۶m۶m�?�$I�$I�?      �?                      �?              �?      �?              �?        ��N��N�?�؉�؉�?�������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?��D�o-�?��n���?�?�������?%I�$I��?�m۶m��?��FS�׾?�!�%�?�$I�$I�?n۶m۶�?F]t�E�?/�袋.�?�$I�$I�?۶m۶m�?�q�q�?��8��8�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�q�q�?9��8���?(�����?�5��P�?              �?      �?              �?      �?      �?                      �?�{a���?5�rO#,�?۶m۶m�?�$I�$I�?              �?      �?      �?333333�?�������?      �?      �?              �?      �?        �������?UUUUUU�?              �?      �?                      �?�?�������?�$I�$I�?n۶m۶�?�������?�������?      �?                      �?              �?      �?        d!Y�B�?��7��M�?              �?l�l��?��I��I�?      �?        p�\��?�я~���?              �?{�G�z�?���Q��?      �?                      �?/�����?h/�����?/�袋.�?F]t�E�?              �?      �?              �?      �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?d!Y�B�?�Mozӛ�?      �?      �?      �?                      �?�����Ң?�������?              �?�������?ffffff�?և���X�?��)x9�?333333�?ffffff�?              �?      �?      �?      �?                      �?              �?      �?        ��`����?�E|���?�H�ls�?��R�O2�?ى�؉��?;�;��?y�5���?Cy�5��?�?�������?              �?      �?              �?        �m۶m��?�$I�$I�?              �?      �?        �������?�������?��2(&�?���|���?��:ڼ�?;ڼOqɀ?�Mozӛ�?d!Y�B�?      �?        �������?UUUUUU�?              �?      �?              �?        �������?�������?Jݗ�V�?�A�Iݷ?�Kh/��?h/�����?UUUUUU�?UUUUUU�?              �?      �?        �������?�?և���X�?9/���?�������?�������?      �?                      �?��.���?F]t�E�?���k(�?(�����?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?        ffffff�?333333�?�������?333333�?      �?                      �?      �?                      �?;�;��?ى�؉��?A�Iݗ��?~ylE�p�?333333�?333333�?              �?�k(���?(�����?      �?        �������?�������?n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?              �?      �?              �?333333�?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?(������?l(�����?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?              �?                      �?^Cy�5�?Q^Cy��?      �?              �?      �?      �?        �$I�$I�?n۶m۶�?UUUUUU�?�������?              �?      �?                      �?      �?      �?�5eMYS�?֔5eMY�?      �?        �A�A�?X|�W|��?              �?�������?�������?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?        ��Moz��?Y�B��?      �?        �������?UUUUUU�?      �?      �?              �?      �?      �?              �?      �?              �?        Y�B��?��Moz��?�������?333333�?              �?      �?        �q�q�?��8��8�?UUUUUU�?UUUUUU�?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK煔h��B�9         �       
             �?2���xA�?J           ��@              U                    �?�l�c!g�?T           ��@               F                    �?z)�J'c�?�            @m@                                  �?�6
����?a             c@                      	          ����?��oh���?/            @R@        ������������������������       �                     ?@                                  �a@�ՙ/�?             E@              	                   d@և���X�?             <@        ������������������������       �                     @        
                           �?      �?             8@                      
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @                                  �_@     ��?             0@        ������������������������       �                      @                                   `@      �?              @        ������������������������       �                     �?                      	          ����?և���X�?             @        ������������������������       �                     @                                  �e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@               #                    �?H�z�G�?2             T@                                  `X@8�Z$���?             :@        ������������������������       �                      @                                  �g@�8��8��?             8@                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               "                    �?���7�?             6@                !                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        $       ;                   �`@X�<ݚ�?!             K@       %       *                   �a@��J�fj�?            �B@        &       )       
             �?r�q��?             @        '       (                   @]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        +       0                    ]@f���M�?             ?@        ,       -                    �?�q�q�?             "@        ������������������������       �                     @        .       /                   �r@      �?             @       ������������������������       �                     @        ������������������������       �                     @        1       :                   hp@�GN�z�?             6@       2       9                    �?�X�<ݺ?
             2@       3       8                    @ףp=
�?             $@       4       7                   �c@      �?              @        5       6                    _@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        <       E                    �Q@@�0�!��?             1@       =       >       
             �?      �?             0@        ������������������������       �                     �?        ?       @                    @O@��S�ۿ?
             .@       ������������������������       �                      @        A       B       	          @33�?؇���X�?             @        ������������������������       �                     @        C       D                    d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        G       N                    �?�>����?.            @T@        H       I                     L@      �?             (@        ������������������������       �                     �?        J       K                   �a@"pc�
�?             &@        ������������������������       �                      @        L       M                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        O       T                   �q@�nkK�?'            @Q@       P       Q                    �?г�wY;�?&             Q@       ������������������������       �                    �I@        R       S                     F@�t����?             1@        ������������������������       �                      @        ������������������������       �        
             .@        ������������������������       �                     �?        V       �                   `f@�ma�H��?�             s@       W       `                   �[@���F6��?�            �r@        X       Y                    Y@�q�q�?             2@        ������������������������       �                     @        Z       [                   �`@��
ц��?             *@        ������������������������       �                     @        \       ]                    l@�<ݚ�?             "@        ������������������������       �                     �?        ^       _       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        a       |                   �b@ rpa�?�            pq@       b       u       	          ����?XB���?�            Pp@        c       t                   0a@�8��8��?<             X@       d       k                    l@�����H�?.             R@       e       f                   pi@�O4R���?            �J@       ������������������������       �                     C@        g       j                   �X@��S�ۿ?             .@        h       i       	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        l       s                    �O@p�ݯ��?             3@       m       n                   �l@�t����?             1@        ������������������������       �                     @        o       p                    �?؇���X�?             ,@       ������������������������       �        
             &@        q       r                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     8@        v       {                    �?��ϩ}��?m            �d@        w       x                   `a@�C��2(�?	             &@       ������������������������       �                      @        y       z                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        d            @c@        }       ~       	          433�?�q�q�?             2@        ������������������������       �                     @               �                    @F@z�G�z�?	             .@       �       �                    �?      �?              @        ������������������������       �                     @        �       �       	          033@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        �       �                   `c@=87��?�            �w@        �       �                    �?      �?              F@       �       �                    �?�q�q�?             8@       �       �                     P@�	j*D�?	             *@       �       �                    �?      �?              @       �       �                   �_@      �?             @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                     L@      �?             @       �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    c@�C��2(�?             &@       ������������������������       �                     "@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?P���Q�?             4@       �       �                   c@�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?>�1�K�?�            �t@       �       �                   �s@�����?�            �q@       �       �                   0h@��u5�?�            �p@       �       �                   �b@`!?��?�            �p@        �       �                   �a@0�z��?�?T             _@       ������������������������       �        9             T@        �       �                   �n@���7�?             F@       ������������������������       �                     9@        �       �                    _@�KM�]�?
             3@        �       �                   �a@      �?              @        ������������������������       �                     �?        �       �       	          ����?؇���X�?             @        ������������������������       �                     @        �       �                    �L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        �       �       	          ���@�5?,R�?W             b@       �       �                    @L@,�d�vK�?V            �a@       �       �                    �?�8���?F             ]@        �       �                   �b@��s����?             5@       �       �                   �e@�KM�]�?             3@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                      @        �       �                    @G@ r���?8            �W@       ������������������������       �        #            �O@        �       �                   �n@      �?             @@        �       �                   �c@�r����?
             .@        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     1@        �       �                   �d@���B���?             :@       �       �                   �p@�n_Y�K�?
             *@       �       �                    @M@�q�q�?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �i@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   @c@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                      @        �       �                   u@ҳ�wY;�?             1@        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    �?�[�IJ�?            �G@       �       �       	          ����?"pc�
�?            �@@        �       �                   �`@�eP*L��?	             &@       �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �K@r�q��?             @        ������������������������       �                     @        �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        ������������������������       �        	             ,@        �t�bh�h)h,K ��h.��R�(KK�KK��hb�Bp  �W���?8T��p�?�d�+H�?�5�m�?�)��)��?7k�6k��?�D�D��?�]�]�?����?ȏ?~��?              �?�a�a�?�<��<��?�$I�$I�?۶m۶m�?      �?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?                      �?ffffff�?333333�?;�;��?;�;��?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?�.�袋�?F]t�E�?UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?r�q��?�"�u�)�?к����?UUUUUU�?�������?      �?      �?              �?      �?                      �?��RJ)��?��Zk���?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �袋.��?]t�E�?��8��8�?�q�q�?�������?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?                      �?�������?ZZZZZZ�?      �?      �?      �?        �?�������?              �?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        h/�����?�Kh/��?      �?      �?      �?        F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?        d!Y�B�?�Mozӛ�?�?�?              �?�?<<<<<<�?      �?                      �?      �?        k�k��?��G��G�?ogH���?�v�ļ�?UUUUUU�?UUUUUU�?              �?�؉�؉�?�;�;�?      �?        �q�q�?9��8���?      �?              �?      �?      �?                      �?�n�ᆫ?Hy�G�?�{a���?GX�i���?UUUUUU�?UUUUUU�?�q�q�?�q�q�?�x+�R�?:�&oe�?              �?�?�������?�������?�������?              �?      �?                      �?Cy�5��?^Cy�5�?�������?�������?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�0��x?Ο��Y��?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?      �?              �?      �?      �?      �?                      �?              �?r�q��?�q�q�?      �?                      �?��N>:��?����?      �?      �?�������?�������?vb'vb'�?;�;��?      �?      �?      �?      �?      �?      �?              �?      �?                      �?      �?      �?      �?      �?      �?                      �?      �?              �?        F]t�E�?]t�E�?              �?      �?      �?              �?      �?        �������?ffffff�?�?�?              �?      �?                      �?�w��5�?�!�c)�?�fӍo�?_�d���?�ߦ5��?��:W�?A��~5�?�1���?|���{�?�B!��?      �?        �.�袋�?F]t�E�?      �?        �k(���?(�����?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        �q�q�?�q�q�?��9�h��?�z2~�Գ?j��FX�?a���{�?z��y���?�a�a�?�k(���?(�����?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?9�{n�S�?�X�0Ҏ�?      �?              �?      �?�������?�?              �?      �?              �?        ��؉���?ى�؉��?;�;��?ى�؉��?UUUUUU�?UUUUUU�?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?      �?                      �?              �?�������?�������?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?        m�w6�;�?���
b�?F]t�E�?/�袋.�?t�E]t�?]t�E�?�������?�������?      �?                      �?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���HhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@C         �       	          033�?SH7�j�?C           ��@              I                    �?��<1G�?@           �@                                  �i@~	~���?{            �h@                      
             �?��a�n`�?:            @W@                     	            �?��?^�k�?)            �Q@       ������������������������       �                     L@               
                   �a@؇���X�?
             ,@               	                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?8����?             7@                                 �_@��
ц��?             *@                                  @O@      �?              @                                  �?؇���X�?             @                                   �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@                                   �[@Lu���}�?A            �Y@                                  @b@�q�q�?             8@                                  �?��s����?             5@                     
             �?�X�<ݺ?	             2@                                   Y@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     @        !       H                     P@H���I�?5            �S@       "       3       
             �?��x�5��?1            @Q@        #       ,                    �?�t����?             A@        $       %                   �^@�q�q�?             "@        ������������������������       �                     �?        &       +                    f@      �?              @       '       (                   �`@؇���X�?             @        ������������������������       �                     @        )       *                   pb@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        -       .       	          433�?`2U0*��?             9@       ������������������������       �                     2@        /       2                   �a@؇���X�?             @        0       1                     L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        4       E                    @M@">�֕�?            �A@       5       6                    �C@>���Rp�?             =@        ������������������������       �                     @        7       D                    @J@�q�q�?             8@       8       9                   �a@p�ݯ��?             3@        ������������������������       �                     @        :       C                    �?��
ц��?
             *@       ;       >                   �d@�eP*L��?	             &@        <       =                   �_@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       @                   pf@r�q��?             @        ������������������������       �                     @        A       B                    a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        F       G                   �_@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        J       i                    �?r�'�Z�?�            �s@        K       ^                    c@�˹�m��?^             c@       L       U       
             �?��.N"Ҭ?T            @a@        M       N                    T@z�G�z�?
             .@        ������������������������       �                     �?        O       P                   `m@؇���X�?	             ,@        ������������������������       �                     @        Q       R                   �b@����X�?             @        ������������������������       �                     �?        S       T                    @L@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        V       ]                    _@ �|ك�?J            �^@        W       X                    �?��v$���?%            �N@        ������������������������       �                     :@        Y       Z       	            �?��?^�k�?            �A@       ������������������������       �                     @@        [       \       	          pff�?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        %             O@        _       `                    �?և���X�?
             ,@        ������������������������       �                     @        a       b       
             �?���!pc�?             &@        ������������������������       �                     @        c       d                    �J@և���X�?             @        ������������������������       �                      @        e       f                   �c@z�G�z�?             @        ������������������������       �                      @        g       h                   `r@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        j       }       
             �?ʔ�k��?g            �d@        k       r                    �?~���L0�?            �H@        l       m       	          ���ٿ����X�?	             ,@        ������������������������       �                     �?        n       o                    _@�θ�?             *@        ������������������������       �                     @        p       q                    @N@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        s       x                   �d@؇���X�?            �A@       t       u                   �b@ ��WV�?             :@       ������������������������       �                     5@        v       w                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                   @e@X�<ݚ�?             "@        ������������������������       �                     @        {       |                   `g@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ~       �                    @M@,Z0R�?H             ]@              �                   @[@p�C��?7            �V@        �       �       	          `ff�?����X�?             @       �       �                    m@r�q��?             @       ������������������������       �                     @        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        1             U@        �       �                    �? �o_��?             9@       �       �                    �M@�q�q�?             5@        ������������������������       �                     @        �       �                    �?      �?             0@       �       �                    c@@4և���?
             ,@       ������������������������       �                     $@        �       �                   �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   `Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?           Py@       �       �                    Z@�"P��?�            �r@        �       �                    �?      �?             $@       �       �                   �`@      �?              @       �       �                    �M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   {@`�g�ɦ�?�            �q@       �       �                   �a@�Q�p6м?�            �q@       �       �       
             �?�:+�X��?u            �g@       �       �                   P`@x��-�?a            �c@       �       �                    �?4��?�?A             Z@       �       �                    �?؇���X�?0            �Q@        �       �                   �q@��
ц��?             *@        �       �                    `@����X�?             @       �       �                    �P@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�}�+r��?(            �L@        ������������������������       �                     @        �       �                   Xp@ "��u�?"             I@       �       �                    @J@��a�n`�?             ?@        ������������������������       �                     *@        �       �                   �X@r�q��?             2@        ������������������������       �                     �?        �       �                   8p@�t����?             1@       �       �       
             �?      �?             0@        ������������������������       �                     @        �       �                   �\@$�q-�?             *@        �       �                   �k@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     A@        ������������������������       �                     �K@        �       �                   �]@z�G�z�?             >@        ������������������������       �                     &@        �       �       	          033�?�����?             3@        �       �                   �`@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?r�q��?             (@        �       �                    �?�q�q�?             @       �       �       	          ����?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    `P@�eGk�T�?<            �W@       ������������������������       �        3            �T@        �       �       
             �?$�q-�?	             *@       ������������������������       �                     &@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?)O���?J             [@       �       �                   �f@��W3�?/            �Q@        �       �                     O@�����H�?             "@       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@�&�5y�?)             O@       �       �                   @[@���Q �?#            �H@        �       �                    �M@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ��� @^����?             �E@       �       �                   �e@��hJ,�?             A@       �       �                   `q@     ��?             @@       �       �                   �g@ �q�q�?             8@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     4@        �       �       	          `ff�?      �?              @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?�<ݚ�?             "@        ������������������������       �                     �?        �       �                   `d@      �?              @       ������������������������       �                     @        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �       
                   @V������?            �B@       �                         �n@z�G�z�?             >@       �                           �?      �?             4@        �       �                    `@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                    	          `ff�?�r����?             .@                                b@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @              	      	          ����?ףp=
�?             $@                                �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 @Q@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �t�b��      h�h)h,K ��h.��R�(KMKK��hb�B�  ���t��?�~�E)�?b;��$��?;��$���?h�����?�)x9/�?�c�1Ƹ?�s�9��?�A�A�?_�_��?              �?�$I�$I�?۶m۶m�?�$I�$I�?�m۶m��?      �?                      �?              �?8��Moz�?d!Y�B�?�;�;�?�؉�؉�?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?              �?                      �?������?*9/���?�������?�������?z��y���?�a�a�?��8��8�?�q�q�?�������?UUUUUU�?              �?      �?              �?                      �?              �?^-n����?Q�Ȟ���?�Q�g���?0�̵�?�?<<<<<<�?UUUUUU�?UUUUUU�?      �?              �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?              �?        {�G�z�?���Q��?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?_�_��?�A�A�?�i��F�?GX�i���?      �?        �������?�������?^Cy�5�?Cy�5��?      �?        �؉�؉�?�;�;�?t�E]t�?]t�E�?�������?�������?              �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?���Ѭr�?�M �L5�?��P^Cy�?^Cy�5�?�3J���?ہ�v`��?�������?�������?              �?۶m۶m�?�$I�$I�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?                      �?�_��e��?�h
���?.�u�y�?;ڼOqɐ?      �?        _�_��?�A�A�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ۶m۶m�?�$I�$I�?      �?        t�E]t�?F]t�E�?              �?۶m۶m�?�$I�$I�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �בz��?�P�
ŭ�?������?����>4�?�m۶m��?�$I�$I�?              �?ى�؉��?�؉�؉�?      �?        �$I�$I�?۶m۶m�?              �?      �?        �$I�$I�?۶m۶m�?;�;��?O��N���?              �?�������?�������?      �?                      �?�q�q�?r�q��?      �?        UUUUUU�?�������?              �?      �?        �FX�i��?	�=��ܳ?��K��K�?h�h��?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?        
ףp=
�?�Q����?UUUUUU�?UUUUUU�?              �?      �?      �?n۶m۶�?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?              �?      �?              �?        �������?�������?[�R�֯�?��+j�?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?Zƞ�?�T?'���?�ԓ�ۥ�?���@��?�Zk��?�ԟRJ�?��N���?l#֥���?ى�؉��?�N��N��?�$I�$I�?۶m۶m�?�;�;�?�؉�؉�?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?              �?        �������?UUUUUU�?      �?                      �?(�����?�5��P�?              �?���Q��?�G�z�?�c�1Ƹ?�s�9��?              �?UUUUUU�?�������?      �?        �?<<<<<<�?      �?      �?              �?;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?              �?              �?�������?�������?              �?^Cy�5�?Q^Cy��?�$I�$I�?۶m۶m�?              �?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?�X�0Ҏ�?��=�ĩ�?              �?;�;��?�؉�؉�?              �?      �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        9��8���?��8��8�?p�z2~��? �
���?�q�q�?�q�q�?              �?      �?      �?              �?      �?        :�s�9�?�1�c��?9/����?����>4�?UUUUUU�?�������?      �?                      �?�qG��?w�qG��?KKKKKK�?�������?      �?      �?�������?UUUUUU�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?                      �?�q�q�?9��8���?      �?              �?      �?              �?      �?      �?      �?                      �?      �?        o0E>��?�g�`�|�?�������?�������?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?�?�������?�������?�������?              �?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�m۶m��?�$I�$I�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���KhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@A         �                    �?�J���?K           ��@              Y       
             �?�r�����?j           ��@                                  `\@��qqY�?�            �i@               	                    �?������?            �D@                                 �Q@г�wY;�?             A@                                   a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @@        
                           �?؇���X�?             @                                 �]@      �?             @                                  `X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                       	          833�?f`�>�l�?o            �d@                                  pe@"pc�
�?&            �K@                     
             �?8��8���?"             H@        ������������������������       �                     �?                                   �?dP-���?!            �G@       ������������������������       �                     7@                                   �?r�q��?             8@                                  @      �?	             0@                                  �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                  �k@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        !       L                    �?hb�Iy��?I            @[@       "       G                   r@��j���?7            �T@       #       D                    @�萻/#�?/            �P@       $       +                    _@П[;U��?*             M@        %       (                    �?�θ�?             *@       &       '                   @]@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        )       *                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ,       C                   q@�ݏ^���?"            �F@       -       <       	          `ff�?D^��#��?            �D@       .       5                   @l@�c�Α�?             =@        /       0       	          ����?؇���X�?             ,@       ������������������������       �                      @        1       4                   �a@�q�q�?             @       2       3                    �D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        6       7                   �l@���Q��?             .@        ������������������������       �                     @        8       9                   @[@"pc�
�?
             &@        ������������������������       �                     �?        :       ;                   0a@ףp=
�?	             $@       ������������������������       �                     "@        ������������������������       �                     �?        =       B       	          `ff@�8��8��?             (@       >       A                   �`@      �?              @        ?       @                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        E       F                   �a@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        H       K                    �?      �?             0@       I       J                    b@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        M       N                    �?�	j*D�?             :@        ������������������������       �                     &@        O       T                    @L@��S���?             .@        P       Q                   �`@r�q��?             @       ������������������������       �                     @        R       S                   f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        U       V                    �N@�q�q�?             "@        ������������������������       �                     @        W       X                   p@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        Z       �       	          ���@�(SD�?�            Pv@       [       j                   `_@�H�i�?�            �u@        \       c                   �S@�θ�?!             J@        ]       b                   a@�θ�?             *@       ^       _                    [@      �?             @        ������������������������       �                      @        `       a       	          ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        d       i       	             �?�7��?            �C@       e       f                   �^@@-�_ .�?            �B@       ������������������������       �                    �@@        g       h                   @m@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        k       �                     L@�C��2(�?�            �r@       l       q                   �e@���Rp�?�             m@        m       p                   @e@r�q��?             2@       n       o                    @I@      �?             0@       ������������������������       �        
             .@        ������������������������       �                     �?        ������������������������       �                      @        r       �                   �b@ 5x ��?�            �j@       s       t                    �F@ %$��ݞ?}            �h@        ������������������������       �        ;            @W@        u       �                   �_@ f^8���?B            �Y@        v       y                    �?��S�ۿ?            �F@        w       x                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        z       {                   �b@ �#�Ѵ�?            �E@       ������������������������       �                     <@        |       }                    �?�r����?             .@        ������������������������       �                     @        ~       �                   �^@      �?              @              �                    c@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        $             M@        �       �                    �?r�q��?	             2@        ������������������������       �                     $@        �       �                    �E@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �_@
��[��?'            @P@        �       �                   0c@����X�?             ,@       �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    s@>a�����?            �I@       �       �                    b@��p\�?            �D@       ������������������������       �                     =@        �       �       	          ����?      �?	             (@        �       �                    e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             $@       �       �                   �b@r�q��?             @       �       �                   0b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �c@r�,����?�            @v@       �       �                    �?�����	�?�            @u@        �       �       
             �?���Q��?            �A@       �       �                   xt@�4�����?             ?@       �       �                    �?�q�q�?             8@       �       �                   pb@      �?             4@       �       �                   �g@�r����?
             .@        ������������������������       �                     �?        �       �       	          433�?@4և���?	             ,@        �       �       	          ����?r�q��?             @        ������������������������       �                     @        �       �                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `c@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    w@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   i@(��y@[�?�            s@        �       �                   pb@���>4ֵ?G             \@       �       �                    �?�(�Tw�?2            �S@       ������������������������       �        (            �O@        �       �                    �?��S�ۿ?
             .@        �       �                    I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     *@        �       �                     F@�t����?             A@        ������������������������       �                     �?        �       �                   �_@�C��2(�?            �@@       ������������������������       �                     8@        �       �                   �`@�q�q�?             "@        ������������������������       �                      @        �       �       	             �?؇���X�?             @        ������������������������       �                     @        �       �                   �g@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �R@��5�W�?}             h@       �       �                    �K@\�ih�<�?|            �g@        �       �                   0n@�:�]��?>            �Y@        �       �                   �m@x�����?            �C@       �       �       	          ����?>A�F<�?             C@        �       �                    �?�����?             3@       �       �       
             �?���Q��?
             .@       �       �       	             �?�	j*D�?             *@        ������������������������       �                      @        �       �       	             �?z�G�z�?             @        ������������������������       �                      @        �       �       	          ����?�q�q�?             @       �       �                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �F@�}�+r��?             3@        �       �       	             @      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �        $            �O@        �       �                   �\@�������?>             V@        �       �                   @l@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?p#�����?8            �S@        �       �                    �L@8����?             7@        �       �                    �?�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �`@@�0�!��?             1@       �       �                    �?��S�ۿ?             .@       ������������������������       �        
             &@        �       �                    ]@      �?             @       �       �                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?@4և���?&             L@       �       �                   �b@��-�=��?            �C@       ������������������������       �                    �A@        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     @        �                          �?      �?	             0@       �             	             �?؇���X�?             ,@       �                          �?$�q-�?             *@                                 �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��hb�BP  T��p��?Vr9�ǎ�?&F�����?�s�6db�?�֤lM��?���Iٚ�?������?p>�cp�?�?�?      �?      �?      �?                      �?              �?�$I�$I�?۶m۶m�?      �?      �?      �?      �?      �?                      �?              �?              �?�+Q���?%jW�v%�?F]t�E�?/�袋.�?�������?�������?      �?        W�+�ɵ?�����F�?              �?UUUUUU�?�������?      �?      �?      �?      �?      �?                      �?              �?              �?�m۶m��?�$I�$I�?      �?                      �?�߅���?��A��.�?�e�@	o�?o4u~�!�?ï�Dz��?z�rv��?�{a���?��=���?ى�؉��?�؉�؉�?/�袋.�?F]t�E�?              �?      �?              �?      �?              �?      �?        ��I��I�?�[�[�?,Q��+�?�]�ڕ��?5�rO#,�?�{a���?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?333333�?�������?              �?/�袋.�?F]t�E�?              �?�������?�������?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?                      �?              �?              �?              �?9��8���?�q�q�?              �?      �?              �?      �?�m۶m��?�$I�$I�?      �?                      �?      �?        ;�;��?vb'vb'�?              �?�?�������?�������?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?\��[���?��ِ���?�kQŏl�?`�tՁ��?ى�؉��?�؉�؉�?�؉�؉�?ى�؉��?      �?      �?      �?              �?      �?      �?                      �?              �?��[��[�?�A�A�?S�n0E�?к����?      �?              �?      �?      �?                      �?      �?        ]t�E�?F]t�E�?O#,�4��?	�=��ܣ?�������?UUUUUU�?      �?      �?      �?                      �?              �?7��XQ�?�@�Ե�?������?և���X�?      �?        H%�e�?��VCӝ?�������?�?      �?      �?              �?      �?        �/����?�}A_Ч?      �?        �������?�?      �?              �?      �?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?        7r#7r#�?�����?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?�������?�?�]�ڕ��?��+Q��?      �?              �?      �?      �?      �?              �?      �?              �?              �?      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?                      �?Y�JV���?�MmjS��?�?{{{{{{�?�������?333333�?��RJ)��?���Zk��?�������?UUUUUU�?      �?      �?�?�������?      �?        �$I�$I�?n۶m۶�?UUUUUU�?�������?              �?      �?      �?      �?                      �?              �?333333�?�������?      �?                      �?              �?�m۶m��?�$I�$I�?      �?                      �?      �?        dٍ���?�D�n�?�m۶mۦ?%I�$I��?�A�A�?p��o���?              �?�?�������?      �?      �?              �?      �?                      �?�?<<<<<<�?      �?        F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?m.j�;�?e�x�1�?Ai�
��?�%N���?�?}}}}}}�?�A�A�?��o��o�?Cy�5��?������?^Cy�5�?Q^Cy��?�������?333333�?;�;��?vb'vb'�?              �?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?                      �?(�����?�5��P�?      �?      �?              �?      �?                      �?      �?                      �?/�袋.�?t�E]t�?9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �#{���?7a~W��?8��Moz�?d!Y�B�?UUUUUU�?UUUUUU�?      �?                      �?�������?ZZZZZZ�?�?�������?              �?      �?      �?      �?      �?              �?      �?                      �?      �?        �$I�$I�?n۶m۶�?�A�A�?}˷|˷�?              �?      �?                      �?      �?              �?      �?۶m۶m�?�$I�$I�?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ,J�zhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK兔h��B@9         �                   �c@�HK��x�?7           ��@              _                    �?r�����?�           �@              $                    �?�M���4�?�            �u@                      
             �?P�?�+��?\            �b@              
                    @L@���c���?>             Z@                                  xp@@�E�x�?            �H@       ������������������������       �                     B@               	                    �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@                                  `]@x��}�?"            �K@                      
             �?@4և���?             <@        ������������������������       �                      @        ������������������������       �                     :@                                  �a@�5��?             ;@                                 `o@     ��?             0@                                  �?r�q��?             (@       ������������������������       �                     $@        ������������������������       �                      @                                   `P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@                                   �?�7����?            �G@        ������������������������       �                     @                      	          ����?��i#[�?             E@       ������������������������       �                     7@               !                    V@�����?             3@                      	             �?d}h���?             ,@                                 �a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        "       #                   �a@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        %       B       
             �?�<ݚ�?{            �h@        &       ?                    �?D�n�3�?$            �L@       '       (                   �[@��6���?             E@        ������������������������       �                     @        )       8                    @�e����?            �C@       *       /                    [@������?             ;@        +       .                   �X@      �?             @        ,       -                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        0       1                    �?�㙢�c�?             7@        ������������������������       �                     "@        2       7                    @L@����X�?
             ,@       3       6                    �?X�<ݚ�?             "@       4       5                     H@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        9       >       	          ���@      �?             (@       :       ;                    �?"pc�
�?             &@        ������������������������       �                     �?        <       =                   �b@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     �?        @       A                    �?��S�ۿ?
             .@        ������������������������       �                     �?        ������������������������       �        	             ,@        C       T                    �?d���i�?W            �a@       D       M                   �_@P�2E��?N            @`@        E       H                    �?     ��?             @@        F       G                   �n@      �?             @       ������������������������       �                     @        ������������������������       �                     @        I       L                   �S@$�q-�?             :@        J       K                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        N       S                   @[@@uvI��?>            �X@        O       P                    �F@؇���X�?             @       ������������������������       �                     @        Q       R                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        9            �V@        U       Z                   �a@�eP*L��?	             &@       V       Y                    `@r�q��?             @        W       X                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        [       \                    �?z�G�z�?             @        ������������������������       �                      @        ]       ^                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        `       q                   �j@�D�d@6�?�            Pv@        a       b                   �_@ �#�Ѵ�?h            �e@       ������������������������       �        B             [@        c       p                    �?      �?&             P@       d       o                   �f@:	��ʵ�?            �F@        e       n       	             @D�n�3�?             3@       f       m                    �N@և���X�?
             ,@       g       l                   �a@���!pc�?             &@       h       i                    �?�����H�?             "@       ������������������������       �                     @        j       k                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �                     3@        r       {                    �?zI�^�p�?n             g@        s       z       
             �?X�<ݚ�?             2@       t       u                    n@      �?             0@        ������������������������       �                     @        v       w                    �?�q�q�?
             (@       ������������������������       �                     @        x       y                     L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        |       �       	          ����?3��e��?_            �d@        }       �                    �?�BbΊ�?!             M@       ~       �                   @\@��E�B��?            �G@               �                   @b@�n_Y�K�?             *@       �       �                    �?����X�?             @        �       �                   �k@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?г�wY;�?             A@       ������������������������       �                     8@        �       �                    �?ףp=
�?             $@       ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       
             �?"pc�
�?             &@       �       �                    �?�<ݚ�?             "@       �       �       	          `ff�?      �?              @        ������������������������       �                     @        �       �                   o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0c@бK/eh�?>            @[@       �       �                    _@@3����?=             [@        �       �                    �? 	��p�?             =@       ������������������������       �                     8@        �       �       
             �?���Q��?             @        ������������������������       �                      @        �       �                     M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        .            �S@        ������������������������       �                     �?        �       �                    @L@v�XԖ�?�            �j@       �       �                   �c@B�xX�?j            `d@        �       �                   �e@      �?              @        ������������������������       �                     @        �       �                    �?      �?             @       �       �                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @J@�1)Vz��?e            `c@       �       �                    �?��F���?X            �`@        �       �                    �I@X�<ݚ�?             ;@       �       �                    �?�LQ�1	�?             7@        ������������������������       �                     "@        �       �                   �f@և���X�?             ,@       �       �                   �\@���!pc�?
             &@        ������������������������       �                     @        �       �                    �?      �?              @       �       �                   �b@      �?             @       �       �                    @G@���Q��?             @       �       �                     D@      �?             @        �       �                    �B@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?����?E            �Z@        �       �       	          ���@�q�q�?             8@       �       �                    ]@�㙢�c�?             7@        �       �                   `\@      �?             @       �       �       
             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �n@�IєX�?             1@       ������������������������       �        	             ,@        �       �                   �d@�q�q�?             @        ������������������������       �                     �?        �       �                   q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        5            �T@        ������������������������       �                     6@        �       �                   �t@Rg��J��?             �H@       �       �                   d@�ՙ/�?             E@        �       �                    �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                    �?���!pc�?            �@@        �       �                    �?؇���X�?	             ,@       �       �                   �`@����X�?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �       
             �?p�ݯ��?             3@        ������������������������       �                     $@        �       �                    �N@�<ݚ�?             "@       �       �                     M@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�BP  �T8q���?��cG��?�Zc�7��?�RNd6�?F �]���?s�7D���?�`Q�(X�?�Oק���?�;�;�?;�;��?9/���?և���X�?              �?;�;��?�؉�؉�?      �?                      �?A��)A�?pX���o�?�$I�$I�?n۶m۶�?      �?                      �?/�����?h/�����?      �?      �?�������?UUUUUU�?      �?                      �?      �?      �?              �?      �?                      �?]AL� &�?G}g����?      �?        �a�a�?�<��<��?      �?        ^Cy�5�?Q^Cy��?۶m۶m�?I�$I�$�?      �?      �?              �?      �?                      �?333333�?�������?      �?                      �?9��8���?�q�q�?(������?l(�����?b�a��?=��<���?              �?�-��-��?�A�A�?B{	�%��?{	�%���?      �?      �?      �?      �?              �?      �?                      �?�7��Mo�?d!Y�B�?      �?        �m۶m��?�$I�$I�?r�q��?�q�q�?�������?UUUUUU�?      �?                      �?              �?      �?              �?      �?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?              �?        �?�������?      �?                      �?v{�e��?P$�Ҽ��?_�^��?z�z��?      �?      �?      �?      �?      �?                      �?�؉�؉�?;�;��?333333�?�������?              �?      �?              �?        �Cc}h��?9/���?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?      �?        t�E]t�?]t�E�?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?���й?}��|���?�}A_Ч?�/����?              �?      �?      �?l�l��?��O��O�?(������?l(�����?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?�q�q�?�q�q�?      �?              �?      �?              �?      �?                      �?              �?              �?              �?              �?�5!({_�?���5!(�?r�q��?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?        S&���?6�'���?���=��?�{a��?AL� &W�?�l�w6��?ى�؉��?;�;��?�m۶m��?�$I�$I�?      �?      �?              �?      �?              �?                      �?�?�?              �?�������?�������?              �?      �?      �?      �?                      �?/�袋.�?F]t�E�?9��8���?�q�q�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ��A��.�?��]8��?h/�����?���Kh�?�{a���?������?              �?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        ���s�?��sHM0�?��(��I�?��\w���?      �?      �?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?~\�ǅ}�?=���?��9����?�d\�?r�q��?�q�q�?Nozӛ��?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?t�E]t�?F]t�E�?              �?      �?      �?      �?      �?333333�?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?              �?      �?                      �?��`��}�?�V�9�&�?UUUUUU�?�������?�7��Mo�?d!Y�B�?      �?      �?      �?      �?              �?      �?                      �?�?�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?      �?              �?        ��S�r
�??4և���?�a�a�?�<��<��?9��8���?�q�q�?      �?                      �?t�E]t�?F]t�E�?�$I�$I�?۶m۶m�?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?Cy�5��?^Cy�5�?              �?9��8���?�q�q�?333333�?�������?      �?                      �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ_vhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM	hzh)h,K ��h.��R�(KM	��h��B@B         �                    �?�HK��x�?A           ��@              -                   �`@���$%��?O           ؀@               "       
             �?�����?j             f@                     	          ����?H%u��?A             Y@        ������������������������       �                    �G@                                   �?�T`�[k�?$            �J@                      
             �?�eP*L��?             &@        ������������������������       �                     �?        	                          �a@      �?             $@       
              	          ����?r�q��?             @       ������������������������       �                     @                                  @^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                    Q@؇���X�?             E@                                 8w@��-�=��?            �C@                                 `]@�˹�m��?             C@        ������������������������       �                     2@                      
             �?R���Q�?             4@        ������������������������       �                      @                                    O@�X�<ݺ?
             2@       ������������������������       �                     *@                                  �_@z�G�z�?             @        ������������������������       �                     @                                  0k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                  �N@�q�q�?             @        ������������������������       �                     �?                !                    �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        #       (                   @c@�=A�F�?)             S@        $       '                    �?�E��ӭ�?	             2@       %       &                    �N@�n_Y�K�?             *@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        )       *                   �^@XB���?              M@       ������������������������       �                    �C@        +       ,                   `_@�KM�]�?             3@        ������������������������       �                      @        ������������������������       �        
             1@        .       c       
             �?�S`���?�            �v@        /       D                    �?8�A�0��?H            �[@        0       5                    �?�Gi����?            �B@        1       2                    �?�<ݚ�?             "@        ������������������������       �                     @        3       4                    r@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        6       7                    �?����X�?             <@        ������������������������       �                     @        8       ?       	          ����?�ՙ/�?             5@       9       :                   �_@����X�?	             ,@        ������������������������       �                      @        ;       <                   �b@�q�q�?             @        ������������������������       �                     @        =       >                   p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        @       A                   0b@և���X�?             @        ������������������������       �                     �?        B       C                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        E       b                    �?X~�pX��?0            @R@       F       [                    �?҄��?+            �P@       G       J                    �?�[�IJ�?            �G@        H       I                    �K@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        K       Z                   �f@�xGZ���?            �A@       L       U                   �c@��S���?             >@       M       R                   �`@���Q��?             4@       N       Q       	          ����?8�Z$���?             *@       O       P                   �b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        S       T                    @E@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        V       Y                    @J@z�G�z�?             $@       W       X                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        \       a                    �J@�S����?             3@        ]       `                    @      �?             @       ^       _       	          ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             *@        ������������������������       �                     @        d       �       	          ����?pe7����?�            �o@       e       �                    �L@��Q�Vz�?�            �l@       f       i                   �O@P���Q�?{             i@        g       h                    �?z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        j       u                    �?��s��?v            �g@        k       p                    �?�㙢�c�?             7@        l       m                   �c@և���X�?             @        ������������������������       �                      @        n       o                   0j@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        q       r                   �g@      �?
             0@       ������������������������       �                     ,@        s       t                    �D@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        v                          �f@ d��?f            �d@       w       x                   Hp@ i�*$Ŋ?`             c@       ������������������������       �        M            �^@        y       ~                    �?(;L]n�?             >@       z       }                   �a@`2U0*��?             9@        {       |                    _@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     3@        ������������������������       �                     @        �       �                    �?z�G�z�?             .@        ������������������������       �                     @        �       �                    @D@���!pc�?             &@       �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    k@8^s]e�?             =@        �       �                    @M@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�+e�X�?             9@        �       �                    �M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ףp=
�?             4@       ������������������������       �        
             .@        �       �                     @���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�q�q�?             8@       �       �                    �?@4և���?	             ,@        ������������������������       �                      @        �       �                    �N@�8��8��?             (@       ������������������������       �                     @        �       �                    a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?ףp=
�?             $@       ������������������������       �                      @        �       �       	             @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   0c@�6�7��?�            �w@       �       �                    �J@x�ۈp�?�            `u@        �       �                   Hq@j��>��?R            ``@       �       �                    �?�q�q��?<             X@       �       �                    Z@��T|n�?5            �U@        �       �                   0a@�q�q�?             @        ������������������������       �                     �?        �       �       	             �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       
             �?\���(\�?1             T@       �       �                    �?�����H�?,             R@        �       �                     I@�q�q�?             @       �       �                   �k@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �D@���}<S�?)            @Q@        �       �                    �?      �?             0@       �       �                   �`@�q�q�?             (@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �m@�&=�w��?"            �J@       ������������������������       �                     C@        �       �                    �?�r����?
             .@       ������������������������       �                     &@        �       �                   @X@      �?             @        ������������������������       �                     �?        �       �       
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �p@      �?              @       �       �                   �`@r�q��?             @        ������������������������       �                     @        �       �                    �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �       	          ����?�z�G��?             $@       �       �                   k@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   `^@��?^�k�?            �A@        �       �                    �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     >@        �       �       
             �?Lő����?�            `j@       �       �                   Pr@@-�_ .�?{             g@       �       �                   �X@Ћ����?l            �d@        �       �                    \@R���Q�?             4@        ������������������������       �                     �?        �       �                   �W@�KM�]�?             3@        ������������������������       �                     "@        �       �                   @X@z�G�z�?             $@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @n@@��8��?_             b@       �       �                    �O@@䯦s#�?B            �Z@       ������������������������       �        1            �S@        �       �                   pa@ 7���B�?             ;@       ������������������������       �                     :@        ������������������������       �                     �?        �       �                   pn@�}�+r��?             C@        ������������������������       �                     �?        �       �       	          ����?�?�|�?            �B@        �       �                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �A@        �       �       	          ����?��s����?             5@        �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �R@��S�ۿ?             .@       ������������������������       �        
             ,@        ������������������������       �                     �?        �       �       	          hff�?R�}e�.�?             :@        �       �                     O@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �Q@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        	             1@        �                          �?��+��?            �B@       �                         �s@�+e�X�?             9@       �                         `q@��2(&�?             6@       �             	             �?     ��?
             0@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �                           @K@z�G�z�?             @        ������������������������       �                     @                                  M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 q@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        �t�bh�h)h,K ��h.��R�(KM	KK��hb�B�  �T8q���?��cG��?���s�M�?��87d�?�.�袋�?�袋.��?���Q��?)\���(�?              �?"5�x+��?���!5��?t�E]t�?]t�E�?      �?              �?      �?�������?UUUUUU�?      �?              �?      �?      �?                      �?              �?�$I�$I�?۶m۶m�?�A�A�?}˷|˷�?^Cy�5�?��P^Cy�?              �?333333�?333333�?      �?        �q�q�?��8��8�?              �?�������?�������?              �?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?��k(��?6��P^C�?r�q��?�q�q�?ى�؉��?;�;��?              �?      �?                      �?GX�i���?�{a���?      �?        �k(���?(�����?              �?      �?        ZÁا��?My�N���?/�袋.�?颋.���?o0E>��?#�u�)��?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?      �?        �<��<��?�a�a�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?                      �?�B�
*�?�^�z���?N6�d�M�?�d�M6��?m�w6�;�?���
b�?UUUUUU�?UUUUUU�?              �?      �?        �_�_�?�A�A�?�������?�?333333�?�������?;�;��?;�;��?333333�?�������?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?�������?�������?�q�q�?�q�q�?      �?                      �?      �?              �?        ^Cy�5�?(������?      �?      �?      �?      �?              �?      �?              �?                      �?              �?�����T�?��HX�?��4}PX�?
�[|=�?ffffff�?�������?�������?�������?              �?      �?        q�����?�X�0Ҏ�?�7��Mo�?d!Y�B�?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?              �?      �?      �?              �?      �?      �?                      �?~�z��;�?J���冘?������?(�����z?      �?        �������?�?���Q��?{�G�z�?�������?UUUUUU�?              �?      �?              �?              �?        �������?�������?      �?        F]t�E�?t�E]t�?      �?      �?              �?      �?              �?        |a���?	�=����?      �?      �?      �?                      �?R���Q�?���Q��?�������?�������?      �?                      �?�������?�������?      �?        333333�?�������?              �?      �?        �������?�������?n۶m۶�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        �������?�������?              �?      �?      �?      �?                      �?zq� ��?��]�W�?�A|�?�w�A�?�_�	)y�?����a�?UUUUUU�?�������?�5eMYS�?����)k�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?        �������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        d!Y�B�?ӛ���7�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�x+�R�?tHM0���?              �?�?�������?              �?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ffffff�?333333�?�������?333333�?              �?      �?              �?        �A�A�?_�_��?�������?�������?      �?                      �?              �?���&��?��%�k�?к����?S�n0E�?��+Q��?ԮD�J��?333333�?333333�?      �?        (�����?�k(���?              �?�������?�������?�������?333333�?              �?      �?                      �?UUUUUU�?UUUUUU�?�x+�R�?R����?              �?h/�����?	�%����?              �?      �?        (�����?�5��P�?      �?        к����?*�Y7�"�?      �?      �?      �?                      �?              �?�a�a�?z��y���?      �?      �?              �?      �?        �?�������?              �?      �?        �;�;�?'vb'vb�?9��8���?�q�q�?      �?              �?      �?              �?      �?                      �?*�Y7�"�?�S�n�?���Q��?R���Q�?t�E]t�?��.���?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?      �?                      �?�������?�������?              �?      �?                      �?      �?              �?        �t�bub��-     hhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��xhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM	hzh)h,K ��h.��R�(KM	��h��B@B         �       
             �?���ƒ�?E           ��@              w       	          pff�?�8����?S           ��@                                 �`@��E��)�?�            �t@                      	          033�?�D�e���?:            @U@       ������������������������       �        3             S@                                   �?�<ݚ�?             "@        ������������������������       �                     @               	                    \@      �?             @        ������������������������       �                     �?        
                          @`@�q�q�?             @        ������������������������       �                     �?                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               X                   �b@F9i�g�?�             o@                                  g@vp�*�?|             h@                                   �?p�ݯ��?
             3@                                   @H@�θ�?             *@        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     @                                  �e@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               5                    @L@w@���?r            �e@                                    Z@���Lͩ�?5            �R@                                  �o@      �?             @                                 @m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        !       ,                    �?����Q8�?2            �Q@        "       #                   �]@և���X�?             @        ������������������������       �                     �?        $       %                    �?�q�q�?             @        ������������������������       �                     �?        &       '                   `]@z�G�z�?             @        ������������������������       �                      @        (       )                    �?�q�q�?             @        ������������������������       �                     �?        *       +       	          ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        -       .                    �?     ��?+             P@       ������������������������       �        #            �J@        /       4                    �?�C��2(�?             &@        0       3       	             �?r�q��?             @        1       2                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        6       7       	          ����?r٣����?=            �X@        ������������������������       �                     7@        8       A                    �M@�����?.             S@        9       >                   �`@� �	��?             9@       :       =                    �?      �?	             0@       ;       <                    @M@���Q��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ?       @                   �s@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        B       W                   �p@��x_F-�?            �I@       C       P                    �?����X�?            �A@        D       I                    �?��S���?
             .@        E       F                    �?����X�?             @       ������������������������       �                     @        G       H                    o@      �?             @        ������������������������       �                      @        ������������������������       �                      @        J       K                   �X@      �?              @        ������������������������       �                     �?        L       O                   �`@؇���X�?             @        M       N                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        Q       V                     R@ףp=
�?             4@       R       U       	          @33�?�}�+r��?
             3@        S       T                   p`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �        	             0@        Y       r                   �c@N{�T6�?&            �K@       Z       e                    �?     ��?!             H@        [       \                     E@��.k���?             1@        ������������������������       �                     @        ]       ^                   �^@�n_Y�K�?	             *@        ������������������������       �                     @        _       `                    @G@X�<ݚ�?             "@        ������������������������       �                     @        a       b       	          ����?r�q��?             @       ������������������������       �                     @        c       d                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       m       	          ����?�n`���?             ?@        g       j                   �n@�q�q�?	             .@       h       i                   �_@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @        k       l                   0c@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        n       o                    �?      �?             0@       ������������������������       �                     $@        p       q                   �\@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        s       v                   pl@؇���X�?             @        t       u                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        x       y                   �U@�`��H �?w            �h@        ������������������������       �                     �?        z       {                   �j@�"P��?v            �h@        ������������������������       �        &            �N@        |       �                   `d@��)��g�?P             a@       }       �                    �?HVĮ���?J            �_@        ~                           �?�n_Y�K�?	             *@       ������������������������       �                      @        ������������������������       �                     @        �       �                    @`����x�?A            �\@       �       �                    �?�?�|�??            �[@       �       �                    \@ �ׁsF�?6             Y@        �       �                    `Q@ �q�q�?             8@       ������������������������       �                     4@        �       �                   �p@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        )             S@        �       �                   Pn@"pc�
�?	             &@        �       �                    �?���Q��?             @       �       �                     K@      �?             @        ������������������������       �                     �?        �       �                    �P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �L@���Q��?             $@       �       �                    @      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?0�q=�?�             x@        �       �                    �?�IєX�?D            �Y@        �       �                   xt@��2(&�?             6@       �       �                   `Z@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �        
             2@        �       �                   `u@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                     R@x�G�z�?7             T@       �       �                   �s@pY���D�?6            �S@       ������������������������       �        1            �Q@        �       �                   �`@�<ݚ�?             "@        ������������������������       �                     @        �       �                   @a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @E@"��Q���?�            �q@        �       �                   P`@hP�vCu�?            �D@       �       �                    �?R�}e�.�?             :@       �       �       	          033�?r�q��?             2@       �       �                   `\@��S�ۿ?	             .@        �       �                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    \@      �?              @        ������������������������       �                     @        �       �                    �O@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       	          hff�?���Q��?
             .@        �       �                   e@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    b@      �?              @       �       �                    �?r�q��?             @        �       �                    �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�+$�jP�?�            `n@        �       �                    �D@N{�T6�?"            �K@        ������������������������       �                     $@        �       �                    q@��S���?            �F@       �       �       	          ����?:ɨ��?            �@@       �       �                    \@r�q��?             8@        �       �                   Pa@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �d@ףp=
�?             4@       �       �                    �H@z�G�z�?             $@        ������������������������       �                     �?        �       �                   0c@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    @�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        �       �                   �v@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                    @G@��E�B��?r            �g@        ������������������������       �        /            @T@        �             	          033�?,y�xEE�?C            �Z@       �       �                    �G@fhK�4�?=            �X@        �       �                   �n@      �?              @        �       �       	          ����?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �l@؇���X�?8            �V@       �       �                   Pi@ 	��p�?%             M@       �       �                    d@��?^�k�?            �A@       ������������������������       �                     <@        �       �                   �f@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @�LQ�1	�?             7@       �       �                   �j@���N8�?             5@        �       �                   pj@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             .@        ������������������������       �                      @        �       �                    @J@���!pc�?            �@@        �       �       	          ����?���|���?             &@       �       �                   `a@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    `@�C��2(�?             6@        ������������������������       �                     �?        �                          �?���N8�?             5@       �                           �O@�}�+r��?             3@       ������������������������       �        	             ,@                                 `@z�G�z�?             @        ������������������������       �                     @                                Pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                �g@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM	KK��hb�B�  �j�1N�?�J.g���?�qA��?��o��9�?��/�]�?��t�h�?�???????�?              �?�q�q�?9��8���?              �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �{����?B!��?c�z���?�~����?^Cy�5�?Cy�5��?ى�؉��?�؉�؉�?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ��l���?Ȥx�L�?�K~��?�6�i�?      �?      �?      �?      �?      �?                      �?      �?        ��Vج?O�o�z2�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?     ��?              �?F]t�E�?]t�E�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?|���?>���>�?              �?^Cy�5�?Q^Cy��?�Q����?)\���(�?      �?      �?333333�?�������?      �?                      �?      �?        �q�q�?9��8���?              �?      �?        �?�������?�$I�$I�?�m۶m��?�?�������?�$I�$I�?�m۶m��?              �?      �?      �?              �?      �?              �?      �?              �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?(�����?�5��P�?�������?�������?      �?                      �?              �?      �?                      �?�S�<%��?pX���o�?      �?      �?�?�������?              �?;�;��?ى�؉��?      �?        �q�q�?r�q��?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?        �9�s��?�c�1��?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?�������?333333�?      �?                      �?      �?      �?      �?        �������?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?m�큍޵?R@�O.D�?      �?        [�R�֯�?��+j�?              �?������?/�#EC�?
�B�P(�?_����z�?ى�؉��?;�;��?              �?      �?        Lg1��t�?��,����?к����?*�Y7�"�?{�G�z�?�G�z��?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?F]t�E�?/�袋.�?�������?333333�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?      �?      �?                      �?              �?F�W>��?�ҡ�3�?�?�?��.���?t�E]t�?�5��P�?(�����?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?333333�?a~W��0�?�3���?      �?        9��8���?�q�q�?      �?        333333�?�������?              �?      �?                      �?��V��?��ۥ���?������?��18��?�;�;�?'vb'vb�?UUUUUU�?�������?�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        �������?�������?              �?      �?        333333�?�������?۶m۶m�?�$I�$I�?      �?                      �?      �?      �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        /�����?B{	�%��?�S�<%��?pX���o�?      �?        �?�������?N6�d�M�?e�M6�d�?�������?UUUUUU�?      �?      �?      �?                      �?�������?�������?�������?�������?              �?�q�q�?�q�q�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?        �l�w6��?AL� &W�?      �?        ��/Ċ��?�@�Ե�?,j�J��?P�W
���?      �?      �?�������?�������?              �?      �?              �?        ۶m۶m�?�$I�$I�?������?�{a���?_�_��?�A�A�?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ��Moz��?Y�B��?��y��y�?�a�a�?�������?UUUUUU�?      �?                      �?      �?                      �?F]t�E�?t�E]t�?F]t�E�?]t�E]�?      �?      �?      �?                      �?      �?        ]t�E�?F]t�E�?              �?��y��y�?�a�a�?�5��P�?(�����?      �?        �������?�������?      �?              �?      �?      �?                      �?      �?              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJݳkUhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@?         j                   a@��e�B��?A           ��@               !                   �c@M��-w�?           �z@                                   �?�K�	H�?[             c@                                  I@p�qG�?;             X@              
       
             �?���1j	�?6            �U@                     	          ����?@	tbA@�?+            @Q@       ������������������������       �                     J@               	                    �Q@�IєX�?             1@       ������������������������       �                     0@        ������������������������       �                     �?                                   �?������?             1@                                  �`@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     $@                                    �?�S����?             �L@                                  @K@¦	^_�?             ?@        ������������������������       �                     @                                  `]@8�Z$���?             :@       ������������������������       �        	             0@                      
             �?���Q��?             $@        ������������������������       �                     �?                                  �_@�q�q�?             "@        ������������������������       �                     �?                                   �?      �?              @                                 �]@���Q��?             @        ������������������������       �                     �?                                  �_@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        "       O                   �a@�{����?�            q@       #       8                    �?��e$�?�            `h@        $       7       	          pff�?H�z���?7             T@       %       0                   r@2%ޑ��?0            �Q@       &       /       
             �?\#r��?*            �N@        '       .                    �?և���X�?             ,@       (       )       	             �?���!pc�?	             &@        ������������������������       �                      @        *       +                    �M@�����H�?             "@       ������������������������       �                     @        ,       -                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �G@        1       2                    �?X�<ݚ�?             "@        ������������������������       �                      @        3       6                    @L@����X�?             @       4       5       	             �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        9       J       	          ����?�LQ�1	�?K            �\@        :       =                   �Y@�99lMt�?            �C@        ;       <                   0j@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        >       I       
             �?П[;U��?             =@       ?       F                   0a@8����?             7@       @       C                   @s@�<ݚ�?             2@       A       B                    �O@�C��2(�?
             &@       ������������������������       �        	             $@        ������������������������       �                     �?        D       E                   �t@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        G       H                   `m@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        K       N                   �j@�"w����?1             S@        L       M                    @      �?             0@       ������������������������       �                     .@        ������������������������       �                     �?        ������������������������       �        %             N@        P       e       
             �?���B���?0            �S@       Q       R                   �e@pH����?'            �P@        ������������������������       �                      @        S       b                    @$�q-�?&            @P@       T       Y       
             �?`Jj��?$             O@        U       V                    �?"pc�
�?             &@        ������������������������       �                     @        W       X                     Q@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        Z       a                    �H@`'�J�?            �I@        [       \                    ]@"pc�
�?             &@        ������������������������       �                     @        ]       ^                    �?���Q��?             @        ������������������������       �                     �?        _       `       	             �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     D@        c       d                    �Q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        f       i                   t@���!pc�?	             &@       g       h                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        k       �                    �?6�Է��?4           �~@       l       �                    �?d��U���?�            �w@       m       �       
             �?�mG'v��?�            Ps@        n       }                   �b@Hg����?5            �V@        o       p                   Pa@�������?             A@        ������������������������       �                      @        q       t                    �?     ��?             @@        r       s                   @q@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        u       x       
             �?$�q-�?             :@        v       w                   `r@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        y       z                   0a@ �q�q�?             8@       ������������������������       �                     4@        {       |                     O@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ~       �                   �r@      �?              L@              �                    �?և���X�?            �H@        �       �                    �?      �?
             0@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                     �?        �       �       	             �?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                    @G@4���C�?            �@@        ������������������������       �                     @        �       �                    �?|��?���?             ;@       �       �                    �?j���� �?	             1@        �       �                   pe@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        �       �                    @�q�q�?             @        ������������������������       �                     @        �       �                   n@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�z�G��?             $@        �       �                   �c@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �? �o�b��?�            `k@        �       �                   Pq@:ɨ��?            �@@       �       �       	             @��s����?             5@       �       �                    @G@R���Q�?             4@        �       �                   �c@�q�q�?             "@        ������������������������       �                      @        �       �                    @E@؇���X�?             @        ������������������������       �                     @        �       �                    k@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �                     �?        �       �                    �?      �?             (@        �       �                    �?r�q��?             @        �       �                    `@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    s@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   pf@����D��?u            @g@       �       �       	          ����?���E�?k            �e@       ������������������������       �        a            �c@        �       �                    �?�t����?
             1@        ������������������������       �                     @        �       �                    d@r�q��?             (@       ������������������������       �                     @        �       �                   �g@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �_@r�q��?
             (@        ������������������������       �                     @        �       �                    �?�q�q�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@R_u^|�?)            �Q@        ������������������������       �                      @        �       �                    �?��~R���?$            �O@        ������������������������       �                     ?@        �       �                   �O@     ��?             @@        �       �                    �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �       
             �?�J�4�?             9@        ������������������������       �                     @        �       �                   @c@�<ݚ�?             2@        ������������������������       �                     �?        �       �                   p@@�0�!��?             1@       ������������������������       �                     $@        �       �                    e@և���X�?             @       �       �                   `c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?������?H             \@       �       �                   Pd@�S����?4             S@       �       �                   �V@�θV�?/            @Q@        ������������������������       �                     �?        �       �                    �?l��\��?.             Q@        �       �                     K@������?
             .@        �       �                   �a@և���X�?             @        ������������������������       �                     @        �       �                   �b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?�&=�w��?$            �J@       �       �                    @G@      �?             @@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     :@        ������������������������       �                     5@        �       �       
             �?����X�?             @        ������������������������       �                     �?        �       �                     K@r�q��?             @        �       �                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          `ff�?�E��ӭ�?             B@       �       �       	            �?؇���X�?             <@        ������������������������       �                     ,@        �       �                   �[@����X�?             ,@        ������������������������       �                     @        �       �                   �i@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?      �?              @       ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  �������?�������?�3����?�?NC�?�l�l�?�g�g�?�������?UUUUUU�?qG�wĭ?�;⎸#�?ہ�v`��?�%~F��?              �?�?�?              �?      �?        �?xxxxxx�?�$I�$I�?۶m۶m�?      �?                      �?              �?              �?^Cy�5�?(������?�RJ)���?��Zk���?      �?        ;�;��?;�;��?              �?�������?333333�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?�������?333333�?      �?              �?      �?              �?      �?                      �?              �?�M��M��?Y�Y��?��I��I�?�=۳=��?�������?�������?�������?�A�A�?��:��?XG��).�?�$I�$I�?۶m۶m�?F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �q�q�?r�q��?      �?        �$I�$I�?�m۶m��?UUUUUU�?�������?              �?      �?              �?                      �?Y�B��?��Moz��?�o��o��?5H�4H��?�������?�������?      �?                      �?��=���?�{a���?8��Moz�?d!Y�B�?�q�q�?9��8���?F]t�E�?]t�E�?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?333333�?�������?      �?                      �?      �?        (�����?Cy�5��?      �?      �?              �?      �?                      �?ى�؉��?��؉���?z�rv��?�1���?      �?        ;�;��?�؉�؉�?�B!��?���{��?F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?        �?�������?F]t�E�?/�袋.�?              �?�������?333333�?              �?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?t�E]t�?�q�q�?�q�q�?              �?      �?                      �?:l��F:�?�'�xr��?��%N��?V ��c�?5����?�+�	��?��O��O�?�-؂-��?�������?�������?      �?              �?      �?�������?UUUUUU�?      �?                      �?;�;��?�؉�؉�?      �?      �?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?      �?      �?              �?�������?�������?              �?�q�q�?9��8���?              �?      �?        m��&�l�?'�l��&�?      �?        	�%����?{	�%���?�������?ZZZZZZ�?F]t�E�?t�E]t�?      �?                      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?ffffff�?333333�?�������?              �?      �?                      �?      �?        E�}O��?�a�]�?N6�d�M�?e�M6�d�?z��y���?�a�a�?333333�?333333�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?                      �?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?              �?      �?        P?���O�?X`��?m��֡�?Ȥx�L��?      �?        <<<<<<�?�?      �?        �������?UUUUUU�?      �?        333333�?�������?      �?                      �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?        2~�ԓ��?�@�6�?      �?        �u]�u]�?EQEQ�?              �?      �?      �?�$I�$I�?�m۶m��?              �?      �?        �z�G��?{�G�z�?      �?        9��8���?�q�q�?              �?ZZZZZZ�?�������?      �?        �$I�$I�?۶m۶m�?�������?�������?      �?                      �?              �?n۶m۶�?I�$I�$�?^Cy�5�?(������?�Q�g���?̵s���?      �?        �������?------�?�?wwwwww�?�$I�$I�?۶m۶m�?      �?              �?      �?              �?      �?                      �?�x+�R�?tHM0���?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        �q�q�?r�q��?۶m۶m�?�$I�$I�?      �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?      �?      �?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���UhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK텔h��B@;         �                    �?�s����?C           ��@              S       
             �?\��[Y�?L           ��@                                  �g@�nd����?�             k@                                  �`@�p ��?0            �T@                                  �?��[�p�?            �G@        ������������������������       �                     @                                   �?���H��?             E@       ������������������������       �                     ;@        	                          @c@�q�q�?             .@       
                           @G@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @                                   �? >�֕�?            �A@                                  �Y@����X�?             @        ������������������������       �                     @                                  �`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     <@               ,                   �a@+�M��?W            �`@                                   i@      �?#             N@        ������������������������       �                     @                      	          ����?���y4F�?"            �L@        ������������������������       �                     1@               )                   �`@�z�G��?             D@                                  �?���Q��?             9@                                  `X@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @               (                   ``@�<ݚ�?
             2@               !                   �_@@�0�!��?	             1@       ������������������������       �                      @        "       #       
             �?�q�q�?             "@        ������������������������       �                     @        $       '                    �?      �?             @       %       &                   �\@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        *       +                     @�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        -       L                   Hr@؀�:M�?4            �R@       .       K                     P@*;L]n�?+             N@       /       J                   @q@H(���o�?(            �J@       0       E       	          ���@~���L0�?$            �H@       1       4                   �h@:�&���?            �C@        2       3                   �^@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        5       >                   �`@��hJ,�?             A@       6       9       	          ����?�>����?             ;@        7       8                   �m@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        :       ;                   �d@�nkK�?             7@       ������������������������       �                     2@        <       =                    �F@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ?       B                    �?և���X�?             @       @       A                    @J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        C       D                   n@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        F       I                   �d@z�G�z�?             $@       G       H                    f@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        M       R                    �?؇���X�?	             ,@       N       Q                   y@����X�?             @       O       P                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        T       _                   @E@D�a���?�            `t@        U       ^                    �?����X�?             <@       V       W                    [@      �?
             0@        ������������������������       �                     @        X       [                     N@�n_Y�K�?	             *@        Y       Z                   `\@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        \       ]                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     (@        `       {                    @L@46��e-�?�            �r@       a       z                    �?��*;�?�             n@       b       w                   0h@p)�����?�             k@       c       d                   �a@p ��g�?�            �j@        ������������������������       �        +            �T@        e       f                    �?�1����?V            ``@        ������������������������       �                    �I@        g       p                   �c@\���(\�?9             T@        h       m                   �c@�	j*D�?             :@       i       j                   �m@�GN�z�?             6@       ������������������������       �        	             &@        k       l                   �^@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @        n       o                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        q       v                    �?�X�<ݺ?&             K@        r       s                   pf@�z�G��?             $@       ������������������������       �                     @        t       u                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     F@        x       y                   pn@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        |       �                    �?����S��?$             M@        }       ~                   �l@
;&����?             7@        ������������������������       �                     @               �                   �b@b�2�tk�?             2@        �       �                   �c@z�G�z�?             @        ������������������������       �                      @        �       �                   �s@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   ps@�θ�?             *@       �       �                    �?      �?              @        ������������������������       �                      @        �       �                   8p@r�q��?             @        ������������������������       �                     @        �       �                    @M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @b�h�d.�?            �A@       �       �                    �L@z�G�z�?             >@        ������������������������       �                     �?        �       �                    �O@д>��C�?             =@       �       �                    �?�X�<ݺ?             2@       �       �                    @M@      �?	             0@       �       �                    c@�����H�?             "@        ������������������������       �                     @        �       �                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �       	          ����?���|���?             &@        ������������������������       �                     @        �       �                    �P@      �?              @        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pd@ l{wY|�?�            �w@       �       �       
             �?�t�~U�?�            �v@       �       �                    �J@d��C��?�            `s@        �       �                   �_@�@��3Z�?>            �X@        ������������������������       �                     I@        �       �                   �n@r�qG�?              H@       �       �                   �k@�'�=z��?            �@@       �       �                    g@�q�q�?             8@       �       �       	          ����?      �?	             0@        ������������������������       �                     @        �       �                    �C@r�q��?             (@        ������������������������       �                     �?        �       �                   `U@�C��2(�?             &@        �       �       
             �?z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    @H@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        �       �                   `Z@ �h�7W�?�            �j@        �       �                   ph@�r����?            �F@       ������������������������       �                     :@        �       �       	          ����?�����?             3@        ������������������������       �                     @        �       �                   �`@��
ц��?             *@        �       �                    _@�q�q�?             "@        �       �                   �j@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��AV���?k            �d@       �       �       
             �? ��ʻ��?W             a@        �       �                   �r@$�q-�?             :@       ������������������������       �                     8@        ������������������������       �                      @        ������������������������       �        H            �[@        �       �                    �N@��� ��?             ?@       �       �                   �a@      �?             0@       �       �                    c@�8��8��?	             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �       	              @      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     .@        �       �                    �?���3�E�?(             J@        �       �                   �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �N@      �?$             H@       �       �                   �a@�q�q�?            �@@       �       �                    �?      �?             6@       �       �       	             �?D�n�3�?             3@        ������������������������       �                     @        �       �       	          033�?d}h���?             ,@       �       �                    �?�8��8��?
             (@        �       �                    �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             &@        �       �                   �a@��S�ۿ?	             .@       ������������������������       �                     (@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �       	          ����?����X�?	             ,@       ������������������������       �                     $@        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  ��mQ��?-I׺��?��)��?��ެ'��?�Kh/��?��Kh/�?��+Q��?Q��+Q�?m�w6�;�?�
br1�?      �?        ��y��y�?�0�0�?              �?UUUUUU�?UUUUUU�?F]t�E�?]t�E�?      �?                      �?      �?        �A�A�?��+��+�?�$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?�n�Wc"�?�HT�n�?      �?      �?      �?        (������?6��P^C�?              �?333333�?ffffff�?�������?333333�?۶m۶m�?�$I�$I�?              �?      �?        �q�q�?9��8���?�������?ZZZZZZ�?              �?UUUUUU�?UUUUUU�?              �?      �?      �?�������?333333�?              �?      �?              �?              �?        �?�������?              �?      �?        E>�S��?v�)�Y7�?""""""�?�������?M0��>��?e�Cj���?����>4�?������?�A�A�?�o��o��?333333�?�������?              �?      �?        KKKKKK�?�������?�Kh/��?h/�����?      �?      �?              �?      �?        �Mozӛ�?d!Y�B�?      �?        �������?�������?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?�q�q�?�q�q�?              �?      �?              �?                      �?              �?۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?�������?UUUUUU�?      �?                      �?              �?      �?        �3���?�0�Qġ�?�$I�$I�?�m۶m��?      �?      �?      �?        ى�؉��?;�;��?      �?      �?      �?                      �?�������?�������?      �?                      �?              �?�m�PM��?R��y�Ź?DDDDDD�?�������?/�����?	�%��Ю?�u&`�X�?u����p�?      �?        J�eDP�?����?      �?        �������?�������?vb'vb'�?;�;��?�袋.��?]t�E�?      �?        t�E]t�?]t�E�?              �?      �?              �?      �?              �?      �?        ��8��8�?�q�q�?ffffff�?333333�?      �?              �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        X�i���?O#,�4��?Y�B��?�Mozӛ�?      �?        9��8���?�8��8��?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �؉�؉�?ى�؉��?      �?      �?      �?        UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?;��:���?_�_��?�������?�������?              �?a���{�?|a���?��8��8�?�q�q�?      �?      �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ]t�E]�?F]t�E�?              �?      �?      �?      �?      �?              �?      �?              �?              �?        ���
b�?���F}g�?��ҟ��?O��I�?�,��?mЦ�?����>4�?���S�r�?              �?�������?�������?|��|�?|���?�������?�������?      �?      �?              �?�������?UUUUUU�?              �?]t�E�?F]t�E�?�������?�������?      �?                      �?      �?                      �?9��8���?�q�q�?      �?                      �?              �?"5�x+��?��sHM0�?�?�������?              �?^Cy�5�?Q^Cy��?              �?�؉�؉�?�;�;�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?7Āt,e�?��8���?�?�������?;�;��?�؉�؉�?              �?      �?                      �?�B!��?�{����?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?              �?b'vb'v�?O��N���?      �?      �?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?      �?(������?l(�����?      �?        ۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?UUUUUU�?�������?              �?      �?                      �?      �?              �?                      �?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �m۶m��?�$I�$I�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�SNhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B@=         n       	          ����?��e�B��?X           ��@                                  �?���7b�?9           `}@                                   �?�7���?S             _@                                  �M@���>4ֵ?J             \@                                 �q@`�E���?@            @X@       ������������������������       �        6            �U@                                   �?z�G�z�?
             $@       ������������������������       �                     @        	       
                   �b@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                   �N@z�G�z�?
             .@        ������������������������       �                     @        ������������������������       �                     (@                                  �`@      �?	             (@                                 �b@�q�q�?             "@        ������������������������       �                      @                      
             �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @               e                    �?���ih)�?�            �u@              4       
             �?�b��[��?�            0q@                                  @f@�>4և��?:             U@        ������������������������       �                     ;@                                   �G@�d�����?(            �L@        ������������������������       �        	             .@               /                   �a@X�Cc�?             E@                                 `h@��S���?             >@        ������������������������       �                     @               "       	          ����?�n_Y�K�?             :@                !                   Pc@@4և���?
             ,@       ������������������������       �        	             *@        ������������������������       �                     �?        #       *                   �m@      �?
             (@        $       %       	          ����?      �?             @        ������������������������       �                     �?        &       '                   �`@�q�q�?             @        ������������������������       �                     �?        (       )                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        +       ,                   q@      �?              @       ������������������������       �                     @        -       .                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        0       1                    @�8��8��?	             (@       ������������������������       �                     "@        2       3                   p@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        5       R                    @L@�,�q��?~            �g@       6       K                    �?8����?c            �b@       7       >                    �?`Ӹ����?Z            �`@        8       =                    �?�q�q�?             (@       9       :                   pe@X�<ݚ�?             "@        ������������������������       �                      @        ;       <                   �p@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ?       @                   pl@�-.�1a�?R            �^@       ������������������������       �        +            @P@        A       B                    @G@XB���?'             M@       ������������������������       �                     >@        C       F                    �?@4և���?             <@        D       E                   @o@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        G       H                    �?�nkK�?             7@       ������������������������       �                     2@        I       J                   �n@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        L       Q                    `@d}h���?	             ,@        M       P                    �I@���Q��?             @       N       O                    �E@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        S       \                    �?�D����?             E@        T       [                   �b@b�2�tk�?             2@       U       Z                    `P@�z�G��?             $@       V       W                    �?      �?              @        ������������������������       �                     @        X       Y                     O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ]       d                   �c@      �?             8@       ^       _                   `a@"pc�
�?             6@        ������������������������       �                     (@        `       a                    �L@���Q��?             $@        ������������������������       �                      @        b       c                    r@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        f       g       
             �?����O��?.            �Q@       ������������������������       �                     F@        h       m                    �?�<ݚ�?             ;@        i       j                    ]@      �?              @       ������������������������       �                     @        k       l                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        o       �                    �?����1�?            |@        p       �       	          ��� @7�A��?p             f@       q       �                    �?�'�=z��?X            �`@        r              
             �?      �?             B@       s       |       	             �?և���X�?             5@        t       {                   �c@z�G�z�?             $@       u       v                   @_@�����H�?             "@        ������������������������       �                     @        w       x                   �]@r�q��?             @        ������������������������       �                     @        y       z                     K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        }       ~                    b@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     .@        �       �                    �?�q�Q�?>             X@       �       �                   �p@      �?(             N@       �       �                   �]@�û��|�?              G@        ������������������������       �                     *@        �       �                    o@�eP*L��?            �@@       �       �       
             �?�	j*D�?             :@       �       �       	          033�?և���X�?             ,@       �       �       	          033�?�q�q�?             "@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �K@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        �       �                     L@؇���X�?             ,@        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �M@tk~X��?             B@        �       �       	          ����?b�2�tk�?             2@        �       �       
             �?؇���X�?             @        �       �                    ^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �X@�eP*L��?             &@        ������������������������       �                     @        �       �                    e@      �?              @       �       �                    �?؇���X�?             @        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@        �       �                    @��2(&�?             F@       �       �                    `@�KM�]�?             C@        ������������������������       �                     1@        �       �                    @O@��s����?             5@        ������������������������       �                     &@        �       �                   �`@���Q��?             $@        ������������������������       �                     @        �       �       	          033@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @b@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   �[@���� �?�             q@        �       �                    g@�LQ�1	�?             7@        ������������������������       �                      @        �       �       	          `ff�?��S���?
             .@       �       �                   �m@�q�q�?             (@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��仞�?�             o@       �       �                    �?����9�?�            �h@        �       �       	          ����?�θ�?             :@        �       �       	          ����?X�<ݚ�?             "@        ������������������������       �                     �?        �       �                    �?      �?              @       �       �                    �H@և���X�?             @        ������������������������       �                      @        �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�t����?
             1@        ������������������������       �                     @        �       �                   �`@8�Z$���?             *@       �       �                   �`@�q�q�?             @        ������������������������       �                      @        �       �                    �I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �       	          033�?Ѝܯ0$�?r            �e@       �       �                   �e@@uvI��?@            �X@        �       �                   pb@������?             B@       ������������������������       �                     =@        �       �                    _@؇���X�?             @        ������������������������       �                     @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        -             O@        �       �                    U@��S�ۿ?2            �R@        �       �                    @M@�<ݚ�?             "@       ������������������������       �                     @        �       �       
             �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    s@���7�?+            �P@       �       �                    �J@@3����?$             K@        �       �                     J@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     E@        �       �                   �\@r�q��?             (@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �`@z�G�z�?             I@        ������������������������       �                     :@        �       �                   �l@�q�q�?             8@        �       �                   �X@�θ�?             *@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     &@        �t�b��     h�h)h,K ��h.��R�(KK�KK��hb�BP  �������?�������?��[�`�?��H�>�?)��RJ)�?��Zk���?%I�$I��?�m۶mۦ??��W�?����?      �?        �������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?              �?      �?              �?      �?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?�����?5�� ��?� O	��?־a��?�m۶m��?�$I�$I�?              �?y�5���?Cy�5��?              �?�m۶m��?%I�$I��?�������?�?      �?        ى�؉��?;�;��?�$I�$I�?n۶m۶�?              �?      �?              �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?      �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?                      �?8���ۤ�?W��l�?`��c.�?�y���??�>��?l�l��?UUUUUU�?UUUUUU�?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?                      �?      �?        {����z�?�h
���?      �?        GX�i���?�{a���?      �?        n۶m۶�?�$I�$I�?�������?�������?              �?      �?        �Mozӛ�?d!Y�B�?      �?        �������?�������?              �?      �?        I�$I�$�?۶m۶m�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �0�0�?z��y���?9��8���?�8��8��?ffffff�?333333�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?      �?/�袋.�?F]t�E�?      �?        333333�?�������?              �?      �?      �?      �?                      �?              �?�]�����? �
���?              �?9��8���?�q�q�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        %I�$I��?�m۶m��?t�E]t�?F]t�E�?|���?|��|�?      �?      �?�$I�$I�?۶m۶m�?�������?�������?�q�q�?�q�q�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        ]t�E�?F]t�E�?      �?                      �?      �?        �������?�������?      �?      �?��,d!�?8��Moz�?              �?t�E]t�?]t�E�?vb'vb'�?;�;��?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?              �?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        9��8���?r�q��?9��8���?�8��8��?�$I�$I�?۶m۶m�?      �?      �?              �?      �?                      �?t�E]t�?]t�E�?              �?      �?      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?                      �?              �?t�E]t�?��.���?(�����?�k(���?              �?�a�a�?z��y���?              �?�������?333333�?      �?        �$I�$I�?۶m۶m�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        <<<<<<�?xxxxxx�?d!Y�B�?Nozӛ��?              �?�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?��"NT��?j�;v5,�?�8���߮?v<���?�؉�؉�?ى�؉��?�q�q�?r�q��?      �?              �?      �?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?              �?�?<<<<<<�?              �?;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?�������?�t�g���?9/���?�Cc}h��?�q�q�?�q�q�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?�?�������?�q�q�?9��8���?              �?      �?      �?              �?      �?        F]t�E�?�.�袋�?h/�����?���Kh�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?              �?�������?�������?ى�؉��?�؉�؉�?      �?      �?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ7G\hhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�?         ~                    �?v�����?F           ��@              +                    �H@�܍�`7�?/           �}@                      
             �?���f��?K            �_@                                  �? �q�q�?,             R@                                  �k@�q�q�?             @        ������������������������       �                     @                                   �?�q�q�?             @        ������������������������       �                     �?        	       
                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   ]@����e��?'            �P@                                   �?�nkK�?             7@                                 �e@��S�ۿ?             .@       ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �E@                                  �e@������?             K@                      	          ����?z�G�z�?             $@                                  0e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @               *                    �?��2(&�?             F@                                  �C@�����?             E@        ������������������������       �                      @                                  �[@�t����?             A@                                   �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                '       	            �?��S�ۿ?             >@       !       "                    �?h�����?             <@        ������������������������       �                      @        #       &                    �?P���Q�?
             4@       $       %                    @D@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �                     0@        ������������������������       �                     @        (       )                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ,       a       	          ����?H~4o]�?�            �u@        -       L                   p`@�J�j�?g            �c@       .       1                    �?�q�q�??             X@        /       0                   �]@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        2       E                    �?H��?"�?8             U@       3       >                    �?r�����?#            �J@       4       =                   �q@      �?             D@       5       <                    b@�˹�m��?             C@       6       ;                    �? �Cc}�?             <@       7       8                   �\@�S����?             3@        ������������������������       �                     @        9       :       
             �?z�G�z�?
             .@       ������������������������       �                     (@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     $@        ������������������������       �                      @        ?       B       
             �?�n_Y�K�?             *@       @       A                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        C       D       	             �z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        F       G       	          `ff�?�g�y��?             ?@       ������������������������       �                     6@        H       I                   pf@�����H�?             "@       ������������������������       �                     @        J       K                     N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        M       Z                    �M@�P�*�?(             O@       N       U                   �a@�Gi����?            �B@       O       R       	             �?�C��2(�?             6@       P       Q                    P@�X�<ݺ?             2@        ������������������������       �                     �?        ������������������������       �        
             1@        S       T                    @M@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        V       Y                    �?�r����?
             .@        W       X                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        [       `                   `f@�J�4�?             9@       \       _                   �h@���7�?             6@        ]       ^                   @h@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     @        b       e       	             �?��ɹ?}            �g@        c       d                    �?�S����?             3@        ������������������������       �                     @        ������������������������       �                     0@        f       q       
             �?�|�%T�?o             e@        g       h                   �W@�ݜ�?            �C@        ������������������������       �                     �?        i       n                   �T@�KM�]�?             C@        j       m                    �O@����X�?             @       k       l                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        o       p                    �R@`Jj��?             ?@       ������������������������       �                     =@        ������������������������       �                      @        r       y                   �c@ ����?U            @`@       s       t       	          033@@���a��?J            �\@       ������������������������       �        :            �W@        u       x                   �_@P���Q�?             4@        v       w                   �\@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        z       }                    �?��S�ۿ?             .@        {       |                    �P@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@               �       	             �?��&�B
�?           �{@       �       �                    I@��2(&�?�            @s@        �       �                    �?�g�y��?             ?@        �       �                   @_@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?����X�?             5@       �       �                     Q@      �?
             0@       ������������������������       �        	             ,@        ������������������������       �                      @        �       �                   �a@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   0h@�.����?�            Pq@       �       �                   �`@`���j��?�             q@       �       �                    @L@ ��^og�?r            �f@       �       �       
             �? �Jj�G�?d            �d@        �       �                    @C@؇���X�?             5@        ������������������������       �                      @        �       �                    �?�}�+r��?             3@       ������������������������       �        
             2@        ������������������������       �                     �?        ������������������������       �        X             b@        �       �                   �d@�E��ӭ�?             2@       �       �                    �L@������?             1@        ������������������������       �                     @        �       �                   �W@@4և���?             ,@        �       �       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             (@        ������������������������       �                     �?        �       �       
             �?������?:            �V@        �       �                    b@p�ݯ��?             3@        �       �                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     O@�eP*L��?             &@       �       �       	          433�?      �?              @       �       �                   0e@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    a@ �q�q�?.             R@        �       �                    �?      �?              @       �       �                    �?����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    c@     ��?*             P@       ������������������������       �                     H@        �       �                    �?      �?             0@        ������������������������       �                     �?        ������������������������       �        
             .@        ������������������������       �                     @        �       �                   �b@(옄��?Y            @a@       �       �                    �?X�Cc�?5             U@       �       �                    �P@և���X�?'            �O@       �       �                    @O@      �?              I@       �       �                    �?���Q��?             D@        �       �                    d@���!pc�?             &@       �       �       
             �?z�G�z�?             $@       �       �                   @_@����X�?             @        �       �       	             �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   s@�c�Α�?             =@       �       �                    @F@���B���?             :@        �       �       	              @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    `@�LQ�1	�?             7@        ������������������������       �                     *@        �       �                   �j@�z�G��?	             $@        ������������������������       �                     @        �       �                   �`@      �?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                   xp@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?ףp=
�?             $@       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @\@8�Z$���?             *@        ������������������������       �                     @        �       �       	          ����?����X�?             @        �       �                   �c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �R@؇���X�?             5@       �       �                    �?�}�+r��?             3@        �       �                   �b@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                      @        �       �                   �\@r�q��?$             K@        ������������������������       �                     @        �       �                   Pc@�t����?"            �I@        ������������������������       �                     "@        �       �       	          033�?؇���X�?             E@        �       �                     @���Q��?             @        ������������������������       �                      @        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @B@������?            �B@        ������������������������       �                     �?        �       �                   �c@�8��8��?             B@       �       �                    �? >�֕�?            �A@       ������������������������       �                     8@        �       �                    @"pc�
�?             &@        ������������������������       �                     @        �       �                    �H@      �?             @        ������������������������       �                     �?        �       �       	          ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  t�W���?�7T���?h8�����?�A�I�?v]�u]��?EQEQ�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?|���?�>����?d!Y�B�?�Mozӛ�?�?�������?              �?      �?                      �?              �?B{	�%��?{	�%���?�������?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?��.���?t�E]t�?=��<���?�a�a�?      �?        <<<<<<�?�?      �?      �?              �?      �?        �������?�?�m۶m��?�$I�$I�?      �?        ffffff�?�������?�?�?              �?      �?              �?              �?      �?              �?      �?                      �?+���}��?5�� ��?D�#{��?^-n����?�������?UUUUUU�?      �?      �?      �?                      �?1�0��?�<��<��?�V�9�&�?Dj��V��?      �?      �?^Cy�5�?��P^Cy�?۶m۶m�?%I�$I��?^Cy�5�?(������?              �?�������?�������?              �?      �?                      �?              �?      �?        ى�؉��?;�;��?      �?      �?      �?                      �?�������?�������?              �?      �?        �B!��?��{���?              �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?�Zk����?�RJ)���?o0E>��?#�u�)��?]t�E�?F]t�E�?��8��8�?�q�q�?              �?      �?              �?      �?      �?                      �?�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?{�G�z�?�z�G��?F]t�E�?�.�袋�?�������?�������?              �?      �?                      �?      �?        m�w6�;�?���\AL�?^Cy�5�?(������?      �?                      �?g\�5�?�9J����?�i�i�?\��[���?      �?        (�����?�k(���?�$I�$I�?�m۶m��?      �?      �?      �?                      �?              �?�B!��?���{��?              �?      �?         �����? �����?���ρ?�uI�ø�?              �?�������?ffffff�?�������?�������?      �?                      �?              �?�?�������?      �?      �?      �?                      �?              �?�C��cw�?�p"�?��.���?t�E]t�?��{���?�B!��?�������?�������?              �?      �?        �$I�$I�?�m۶m��?      �?      �?              �?      �?        �������?�������?      �?                      �?�nh��?�ǈ�d�?꫄�YP�?���s2}�?��Z9��?�"Qj�a�?k߰�k�?��)A��?۶m۶m�?�$I�$I�?              �?�5��P�?(�����?      �?                      �?      �?        �q�q�?r�q��?xxxxxx�?�?              �?n۶m۶�?�$I�$I�?      �?      �?              �?      �?              �?                      �?�������?�Q�Q�?Cy�5��?^Cy�5�?      �?      �?      �?                      �?t�E]t�?]t�E�?      �?      �?      �?      �?      �?                      �?              �?      �?        �������?UUUUUU�?      �?      �?�m۶m��?�$I�$I�?              �?      �?              �?             ��?      �?      �?              �?      �?              �?      �?                      �?���,d�?ӛ���7�?�m۶m��?%I�$I��?۶m۶m�?�$I�$I�?      �?      �?�������?333333�?F]t�E�?t�E]t�?�������?�������?�m۶m��?�$I�$I�?333333�?�������?              �?      �?              �?              �?                      �?�{a���?5�rO#,�?ى�؉��?��؉���?UUUUUU�?UUUUUU�?      �?                      �?Y�B��?��Moz��?              �?333333�?ffffff�?              �?      �?      �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?      �?      �?                      �?      �?        ;�;��?;�;��?              �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?�$I�$I�?۶m۶m�?(�����?�5��P�?      �?      �?              �?      �?                      �?      �?        �������?UUUUUU�?              �?<<<<<<�?�?      �?        ۶m۶m�?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ��g�`��?к����?              �?UUUUUU�?UUUUUU�?��+��+�?�A�A�?      �?        /�袋.�?F]t�E�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�[�hG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyK�hzh)h,K ��h.��R�(KK���h��B�?         �       	          033�?�>�Ļ`�??           ��@              E                    �?j�x)��?*           }@               8                    �?��"�y��?y            �g@                     
             �?П[;U��?Z             b@                      	          ����?�j�'�=�?)            �P@                                  �?���7�?             F@               
                     I@���Q��?             @               	                   �b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                    �C@                                   b@�GN�z�?             6@                                  �I@R���Q�?
             4@                                   �?և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        ������������������������       �                      @               /                    �?�6i����?1            �S@              "                   �c@d�;lr�?&            �O@                                 @E@�:�^���?            �F@                                  �X@���Q��?             @        ������������������������       �                      @                                   �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �n@�(\����?             D@       ������������������������       �                     ?@                                   �?�����H�?             "@        ������������������������       �                     �?                !                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     @        #       .                   @c@b�2�tk�?             2@       $       '                    �?     ��?             0@        %       &                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        (       -                   @d@r�q��?             (@        )       *                   �i@�q�q�?             @        ������������������������       �                     �?        +       ,                   d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        0       7                   �d@     ��?             0@       1       4                   �]@��
ц��?	             *@        2       3                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        5       6                    b@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        9       D                   �p@�㙢�c�?             G@       :       ;                   Pj@��p\�?            �D@       ������������������������       �                     <@        <       A                   ``@�θ�?
             *@       =       @                    �J@�����H�?             "@        >       ?                     I@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        B       C                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        F       y                    �?�uA�?�             q@       G       P                   �c@��(�2Y�?�            �k@        H       I       
             �?     ��?             0@       ������������������������       �                     @        J       K                   �]@X�<ݚ�?             "@        ������������������������       �                      @        L       O                   `_@����X�?             @        M       N                    ^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        Q       d       
             �?�b�E�V�?�            �i@        R       [                   �n@X�Cc�?             <@       S       Z                    @O@@�0�!��?             1@       T       U       	          pff�?      �?
             0@        ������������������������       �                     $@        V       Y                    �L@�q�q�?             @       W       X                    �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        \       c                    a@���|���?	             &@       ]       ^                   �a@      �?              @        ������������������������       �                      @        _       b                   �_@�q�q�?             @       `       a                   Xp@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        e       x                   �g@X;��?v            @f@       f       s                    c@@�E��@�?u            �e@       g       p       	             �?@ o����?m            �d@       h       i                   Hp@ A��� �?k            @d@       ������������������������       �        M             ]@        j       o                   0b@��<b�ƥ?             G@        k       l                    �?      �?             0@       ������������������������       �                     "@        m       n                   �p@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     >@        q       r                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        t       u                   pd@ףp=
�?             $@       ������������������������       �                     @        v       w                   �j@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        z       {       	          ���ٿθ	j*�?             J@        ������������������������       �                      @        |       �                   �_@�z�G��?             I@        }       ~                     G@���!pc�?             &@        ������������������������       �                      @               �       
             �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?:�&���?            �C@        �       �                    �?      �?             ,@       �       �                    `P@���|���?             &@       �       �       	          ����?և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     9@        �       �                    �?zW�]�?           P|@       �       �                    �?�U�=���?�            �t@        �       �                   �e@     8�?(             P@       �       �       
             �?�^����?%            �M@        �       �       	          ����?���Q��?             @        ������������������������       �                     �?        �       �                    �?      �?             @       �       �       	          `ff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �       	          ����?h�WH��?!             K@        �       �                   pr@r�q��?
             2@       �       �                    �O@�t����?	             1@       �       �       
             �?      �?             0@       ������������������������       �                     *@        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    `Q@�X�<ݺ?             B@       �       �                    �?��?^�k�?            �A@        �       �                   �`@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     <@        ������������������������       �                     �?        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   @^@�}�+r��?�            �p@        �       �                   `_@ZՏ�m|�?!            �H@        �       �                   �s@ �q�q�?             8@       ������������������������       �                     7@        ������������������������       �                     �?        �       �                    �? �o_��?             9@        ������������������������       �                     @        �       �                    \@�q�q�?             5@       �       �                     M@�eP*L��?             &@       �       �                   ph@�q�q�?             "@        ������������������������       �                      @        �       �       	             @؇���X�?             @        ������������������������       �                     @        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @N@ףp=
�?             $@       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �D@ ��>χ�?~             k@        ������������������������       �                      @        �       �                    @M@�]�h\��?}            �j@       ������������������������       �        L             `@        �       �                    c@`��F:u�?1            �U@       �       �                   pa@��?^�k�?&            �Q@        ������������������������       �                     =@        �       �                    �M@������?            �D@        ������������������������       �                      @        ������������������������       �                    �C@        �       �       
             �?�t����?             1@       ������������������������       �        
             .@        ������������������������       �                      @        �       �                   �e@j�6�<�?N            �^@        �       �       
             �?�LQ�1	�?             7@        ������������������������       �                     @        �       �                    �N@r�q��?             2@       ������������������������       �        
             ,@        �       �                   p`@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?x��#���?>             Y@        �       �                   ``@�>4և��?             <@        �       �                   @c@�q�q�?             (@        �       �                    �K@����X�?             @        ������������������������       �                     �?        �       �                   0l@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             0@        �       �                    @L@*O���?-             R@        �       �                    _@�ʻ����?             A@        ������������������������       �                      @        �       �                   �l@     ��?             @@        �       �                     I@�8��8��?	             (@        �       �       	             �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?
             4@        ������������������������       �                     @        �       �                   @_@�n_Y�K�?             *@        ������������������������       �                     @        �       �                   �l@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �]@>A�F<�?             C@        �       �                    �O@      �?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �M@      �?             @@        �       �                   �_@���!pc�?             &@        ������������������������       �                      @        �       �                   �c@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �       
             �?���N8�?             5@       ������������������������       �                     2@        �       �                   �a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KK�KK��hb�B�  Qm4��?X��;�?�U$^E��?;T�Cu;�?o��2�|�?H���A�?�{a���?��=���?m��&�l�?�&�l���?F]t�E�?�.�袋�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�袋.��?]t�E�?333333�?333333�?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?kq�w��?T:�g *�?��i��i�?�eY�eY�?}�'}�'�?l�l��?�������?333333�?              �?UUUUUU�?UUUUUU�?              �?      �?        333333�?�������?      �?        �q�q�?�q�q�?      �?              �?      �?              �?      �?        �8��8��?9��8���?      �?      �?      �?      �?              �?      �?        �������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?                      �?      �?      �?�؉�؉�?�;�;�?�������?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?        d!Y�B�?�7��Mo�?��+Q��?�]�ڕ��?              �?�؉�؉�?ى�؉��?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?        �H���?ܺ���?�����?*�Y7�"�?      �?      �?              �?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �jch���?��,�?%I�$I��?�m۶m��?ZZZZZZ�?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?F]t�E�?]t�E]�?      �?      �?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�u�{���?�E(B�?ĦҐs�?E'�卑?�?�����?�0�ӈ?,R�n��?�����Hy?      �?        ��7��M�?d!Y�B�?      �?      �?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?              �?      �?      �?                      �?              �?�؉�؉�?�N��N��?              �?ffffff�?333333�?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?      �?        �A�A�?�o��o��?      �?      �?]t�E]�?F]t�E�?۶m۶m�?�$I�$I�?              �?      �?              �?                      �?      �?        YW.���?*>jt���?e�M6�d�?�M6�d��?      �?     ��?W'u_�?u_[4�?�������?333333�?              �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?B{	�%��?��^B{	�?UUUUUU�?�������?�?<<<<<<�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �q�q�?��8��8�?�A�A�?_�_��?�$I�$I�?۶m۶m�?      �?                      �?              �?      �?        �������?�������?      �?                      �?(�����?�5��P�?9/����?�>4և��?UUUUUU�?�������?              �?      �?        �Q����?
ףp=
�?              �?UUUUUU�?UUUUUU�?t�E]t�?]t�E�?UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?      �?              �?      �?      �?                      �?              �?�������?�������?�������?�������?              �?      �?      �?      �?                      �?              �?�@q�8P�?�u�:~�?      �?        ��0�?sy�7�g�?              �?Ȥx�L��?�u�7[��?�A�A�?_�_��?              �?������?p>�cp�?      �?                      �?�?<<<<<<�?              �?      �?        鰑�?yr�'�x�?Y�B��?��Moz��?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?\���(\�?R���Q�?�$I�$I�?�m۶m��?�������?�������?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?      �?                      �?      �?              �?        �q�q�?�q�q�?�������?<<<<<<�?              �?      �?      �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?      �?        �������?333333�?              �?;�;��?ى�؉��?              �?�q�q�?�q�q�?              �?      �?        Cy�5��?������?      �?      �?              �?      �?              �?      �?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?      �?        �a�a�?��y��y�?              �?UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��uhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyM'hzh)h,K ��h.��R�(KM'��h��B�I         �                    �?�HK��x�?@           ��@              ;       	          ����?��s1�?3           p~@                                    �L@�O6o3-�?d            `c@              	       
             �?�d�~V��?C            @X@                                   �?������?             �D@                                   �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �A@        
                          �U@4և����?#             L@        ������������������������       �                      @                                   �?�{��?��?"             K@        ������������������������       �                     ,@                                   �?��Q���?             D@                                  P@      �?             @@                      	          `ffֿz�G�z�?             @        ������������������������       �                      @                                  `[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   ]@PN��T'�?             ;@                                  g@      �?              @        ������������������������       �                      @                                  �[@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     3@                                   �I@      �?              @       ������������������������       �                     @                                  �l@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        !       :                   f@>���Rp�?!             M@       "       9                   �c@d}h���?              L@       #       6                   8r@������?            �F@       $       /                   @a@x�����?            �C@       %       *                   �Y@��hJ,�?             A@        &       )                    �?      �?              @        '       (                   �\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        +       ,       
             �?$�q-�?             :@       ������������������������       �        
             7@        -       .       	          ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        0       5                    @O@���Q��?             @       1       4                    �M@�q�q�?             @       2       3                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        7       8       
             �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                      @        <       �                   Pe@��Lɿ��?�            �t@       =       V                    �?���}<S�?�             t@        >       Q                   pc@� y���?,            �P@       ?       @                   Pl@X�;�^o�?$            �K@       ������������������������       �                     A@        A       D                   �Z@�q�q�?             5@        B       C                   �^@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        E       N                    �?������?             1@       F       K                   `c@d}h���?             ,@       G       H                   �q@�C��2(�?	             &@       ������������������������       �                      @        I       J                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        L       M                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        O       P                     K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        R       S                   pn@�q�q�?             (@        ������������������������       �                     @        T       U                   xu@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        W       X                   �U@��S�ۿ?�            �o@        ������������������������       �                      @        Y       d                    �?���T��?�            �o@        Z       c                    �N@�q�q�?             8@       [       b                   �a@�t����?             1@       \       a                   �d@      �?             $@       ]       `                    `@      �?              @        ^       _       	             �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        e       �                    c@x���a�?�            �l@       f       s                   @^@��~F�<�?x            �h@        g       r                    �?�8��8��?#             H@       h       i                   `_@(N:!���?            �A@       ������������������������       �                     5@        j       m                   �`@����X�?             ,@        k       l                   �j@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        n       q                   �l@�����H�?             "@        o       p                   Pd@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        t                           �?@m����?U            �b@       u       |                   �b@ _�@�Y�?E             ]@       v       {       	          ����?�Ru߬Α?C            �\@        w       z                    �L@      �?              @        x       y       
             �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        ?            �Z@        }       ~                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �@@        �       �                   �r@      �?             @@       �       �                   `c@ ��WV�?             :@        �       �                     L@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     7@        �       �                    �P@      �?             @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?z�G�z�?             $@       �       �                    �?�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @K@�� {�?           �z@       �       �       	          ���@>n�ƌ�?�            p@       �       �                    �?L����?�            �n@       �       �       
             �?(S;�@�?�            �k@        �       �                   @`@���j��?             G@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   Ph@z�G�z�?             D@        �       �                   �]@�q�q�?             "@        ������������������������       �                      @        �       �                   �a@؇���X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   `a@`Jj��?             ?@       �       �                    �?XB���?             =@        ������������������������       �                     &@        �       �                    @G@�X�<ݺ?
             2@       ������������������������       �                     (@        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                    �I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�d���?u            �e@        �       �                     H@      �?             0@       ������������������������       �                     $@        �       �                    �?�q�q�?             @        ������������������������       �                     @        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        �       �                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   @n@�Fǌ��?h            �c@       ������������������������       �        B            �W@        �       �                    �?      �?&             P@       ������������������������       �                     H@        �       �                    �F@      �?             0@        ������������������������       �                     @        �       �                   �n@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                   �`@�5��?             ;@        ������������������������       �                     @        �       �                    �?���N8�?             5@        ������������������������       �                     @        �       �                    d@�t����?	             1@        ������������������������       �                     @        �       �                   �e@�q�q�?             (@        �       �                   �d@z�G�z�?             @        ������������������������       �                     �?        �       �                    @I@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �       	             �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �       
             �?ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        �                         �c@�S����?g            �e@       �             	          ����?�%�E�?Q            `a@       �       �       	          ����?     ��?7             X@       �       �                   �T@l`N���?            �J@        �       �       
             �?��S�ۿ?             .@       ������������������������       �                     &@        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�s��:��?             C@        �       �                   Hs@@4և���?
             ,@       ������������������������       �        	             *@        ������������������������       �                     �?        �       �                   �`@�q�q�?             8@        �       �                    �?�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        �       �       
             �?@4և���?             ,@       ������������������������       �                     @        �       �                    @؇���X�?             @       �       �                    q@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?��V#�?            �E@       �       �                   �l@�������?             >@       �       �                   @b@      �?	             0@       ������������������������       �                     (@        �       �                   `\@      �?             @       �       �                     L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@և���X�?             ,@       ������������������������       �                     @        �       �                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �       	          ����?��
ц��?             *@        ������������������������       �                     �?        �                           O@�q�q�?             (@       �       �                    �?      �?             $@        ������������������������       �                     @        �             
             �?����X�?             @       �                           �?���Q��?             @        ������������������������       �                      @                                pa@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @                    	          `ff�?&^�)b�?            �E@                               @n@�q�q�?             8@             	                   �L@��
ц��?	             *@        ������������������������       �                     @        
                        �`@�<ݚ�?             "@                                 �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@                                 ]@�}�+r��?             3@                    
             �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             0@                                 �e@��R[s�?            �A@                                �?R���Q�?             4@                                 �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 @M@      �?
             0@       ������������������������       �                     &@                                �`@z�G�z�?             @        ������������������������       �                     @                                 �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        !      &      	          ��� @���Q��?             .@       "      %      	             �?      �?             (@       #      $                   l@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM'KK��hb�Bp  �T8q���?��cG��?ޖ�o��?I����?\�ǅ}\�?�=���?�,O"Ӱ�?�i�n�'�?������?p>�cp�?UUUUUU�?UUUUUU�?      �?                      �?              �?%I�$I��?n۶m۶�?              �?���^B{�?/�����?      �?        333333�?�������?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?&���^B�?h/�����?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?      �?              �?      �?      �?                      �?GX�i���?�i��F�?۶m۶m�?I�$I�$�?�?wwwwww�?�A�A�?��o��o�?�������?KKKKKK�?      �?      �?      �?      �?              �?      �?                      �?;�;��?�؉�؉�?              �?UUUUUU�?UUUUUU�?      �?                      �?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        rY1P»?�������?d!Y�B�?ӛ���7�?~5&��?z�rv��?J��yJ�?�־a��?              �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?�?xxxxxx�?۶m۶m�?I�$I�$�?F]t�E�?]t�E�?              �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?        �q�q�?�q�q�?              �?      �?        �?�������?      �?        qК3[�?�R��N�?�������?UUUUUU�?�������?�������?      �?      �?      �?      �?      �?      �?      �?                      �?      �?                      �?              �?              �?��
�[�?�_OE��?&���0�?�;�Y�?UUUUUU�?UUUUUU�?�A�A�?|�W|�W�?              �?�$I�$I�?�m۶m��?333333�?�������?      �?                      �?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�3�=l}�?2�O
��?�{a���?#,�4�r�?p�}��?���#��?      �?      �?      �?      �?      �?                      �?              �?              �?      �?      �?              �?      �?                      �?      �?      �?;�;��?O��N���?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?              �?      �?        �������?�������?�q�q�?�q�q�?      �?                      �?              �?Ն�z��?W�
���?�d�d�d�?�m�m�m�?�Ň+Z_�?S���.�?��oX���?�S�<%ȳ?ozӛ���?!Y�B�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?              �?���{��?�B!��?GX�i���?�{a���?      �?        ��8��8�?�q�q�?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?              �?      �?      �?                      �?�:���C�?Ȥx�L��?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?1���M��?�3���?      �?              �?      �?      �?              �?      �?      �?        �������?�������?              �?      �?        h/�����?/�����?              �?�a�a�?��y��y�?      �?        �������?�������?      �?        �������?�������?�������?�������?              �?      �?      �?              �?      �?        ۶m۶m�?�$I�$I�?      �?                      �?�������?�������?      �?                      �?�:���C�?��2)^�?��\*�?����j�?      �?      �?
�[���?�R���?�?�������?              �?      �?      �?      �?                      �?��k(��?�k(���?n۶m۶�?�$I�$I�?      �?                      �?UUUUUU�?UUUUUU�?ffffff�?333333�?      �?                      �?�$I�$I�?n۶m۶�?              �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?eMYS֔�?6eMYS��?�������?�������?      �?      �?      �?              �?      �?      �?      �?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?        �$I�$I�?۶m۶m�?      �?                      �?�؉�؉�?�;�;�?      �?        �������?�������?      �?      �?              �?�m۶m��?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�}A_��?���/��?�������?�������?�;�;�?�؉�؉�?              �?9��8���?�q�q�?      �?      �?              �?      �?              �?                      �?(�����?�5��P�?UUUUUU�?UUUUUU�?      �?                      �?              �?X|�W|��?PuPu�?333333�?333333�?      �?      �?      �?                      �?      �?      �?      �?        �������?�������?      �?              �?      �?      �?                      �?333333�?�������?      �?      �?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?�t�bub��R      hhubh)��}�(hhhhhNhKhKhG        hh%hNhJjrhG        hNhG        hNhFKhHKhIh)h,K ��h.��R�(KK��hb�C              �?�t�bhUhghPC       ���R�hkKhlhoKh)h,K ��h.��R�(KK��hP�C       �t�bK��R�}�(hKhyMhzh)h,K ��h.��R�(KM��h��B@A         �       
             �?j���� �?;           ��@              Y                    �?���{�?Q           (�@                      	          ����?���X��?�             l@                      
             �?��(�2Y�?1            �R@        ������������������������       �                      @                                  ``@���Hx�?0             R@                                   �?г�wY;�?             A@       ������������������������       �                     9@        	                          `X@�����H�?             "@        
                           �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  �`@�S����?             C@        ������������������������       �                      @                                  �c@�����H�?             B@        ������������������������       �                     0@                                  �d@z�G�z�?             4@                                  �?X�<ݚ�?	             "@        ������������������������       �                     @                                  �c@z�G�z�?             @       ������������������������       �                     @                                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@               B       	          `ff�?Fx$(�?]            �b@              =                    �P@JJ����?;            �W@              "                    ]@�q�q�?7             U@               !                   �X@��S�ۿ?             .@                                  `X@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        #       :                    �?ꮃG��?,            @Q@       $       9                   Xr@�eP*L��?"            �K@       %       ,                    �?JJ����?            �G@        &       +                     L@�E��ӭ�?	             2@        '       (                    �?����X�?             @        ������������������������       �                     @        )       *                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        -       .                    �D@�f7�z�?             =@        ������������������������       �                     @        /       4                    m@`�Q��?             9@       0       1                   �b@@4և���?             ,@       ������������������������       �                     "@        2       3                   �Q@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        5       6       	          ����?���|���?             &@        ������������������������       �                      @        7       8       	          ����?�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ;       <                    �J@����X�?
             ,@        ������������������������       �                     @        ������������������������       �                     $@        >       ?                   �_@ףp=
�?             $@        ������������������������       �                     @        @       A                   @`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        C       D                    �?4և����?"             L@        ������������������������       �                     :@        E       L       
             �?*;L]n�?             >@        F       G                   @]@���!pc�?             &@        ������������������������       �                      @        H       K                    @�����H�?             "@        I       J                   @_@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        M       R                    �?�d�����?             3@       N       Q                   �`@�C��2(�?             &@        O       P                     H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        S       T                    �L@      �?              @        ������������������������       �                     @        U       V                   `b@z�G�z�?             @        ������������������������       �                     @        W       X                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Z       k                    �?Dd�����?�            Pt@        [       `                    �J@����>�?            �B@        \       ]       	          ����?�n_Y�K�?             *@        ������������������������       �                     @        ^       _                    �I@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        a       j                     O@�8��8��?             8@       b       i                     N@�t����?             1@       c       h                    �L@      �?             0@       d       e                    �K@؇���X�?             @        ������������������������       �                     @        f       g                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        l       o                    Z@�8��8��?�             r@        m       n                   0a@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                      @        p                          �[@p��%���?�            @q@        q       t                    �?      �?             8@        r       s                    �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        u       v                   `_@�S����?             3@       ������������������������       �                     $@        w       ~                    �?�q�q�?             "@       x       }                    �?և���X�?             @       y       |                   �k@      �?             @       z       {                    �G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �b@ ,V�ނ�?�            �o@       �       �                    �R@0�M�n�?�             n@       �       �                    �?0�����?�            �m@       �       �                    \@�M����?�            @i@        �       �                   �[@�nkK�?/            @Q@       �       �                   0p@��v$���?*            �N@       ������������������������       �                      G@        �       �                    Z@��S�ۿ?
             .@       ������������������������       �                     (@        �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �       	             @      �?              @       ������������������������       �                     @        �       �                     M@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        Q            �`@        �       �                   �e@�L���?            �B@       �       �                   P`@�IєX�?             A@       �       �                   �_@�t����?
             1@       ������������������������       �                     *@        �       �                    �?      �?             @       �       �                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     1@        �       �                    b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                     M@"pc�
�?             &@       �       �                   �l@ףp=
�?             $@        �       �                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @E@ԛ�c��?�            w@        �       �                    �?�q����?             �J@        �       �                   �X@��H�}�?             9@        ������������������������       �                     @        �       �                    �?���N8�?             5@        �       �                   @b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?r�q��?	             2@       �       �       	          hff�?�r����?             .@       ������������������������       �                     *@        ������������������������       �                      @        �       �                   b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     <@        �       �       	          pff�?��ܾ�"�?�            �s@       �       �                    @L@�|K��2�?�             p@       �       �                    �?�X�<ݺ?�            �h@       �       �                   �f@`�q�0ܴ?}            �g@       �       �                   `\@�g�y��?|            @g@        �       �                   �h@,���i�?            �D@        �       �                    �?      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�FVQ&�?            �@@       ������������������������       �                     0@        �       �                    �?�t����?
             1@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    �H@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    @D@ ���?b             b@        �       �                    �?��?^�k�?            �A@        ������������������������       �                     @        �       �                    �?(;L]n�?             >@        ������������������������       �                      @        �       �                   �b@h�����?             <@       ������������������������       �                     :@        �       �                   Pe@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        K            �[@        ������������������������       �                      @        �       �                    �H@�z�G��?             $@        �       �                   �n@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �a@      �?&             N@        �       �                    @P���Q�?             4@       ������������������������       �                     1@        �       �                    ^@�q�q�?             @        ������������������������       �                     �?        �       �                   ``@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?��Q��?             D@        �       �                   �r@      �?
             0@       �       �                   �_@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �a@      �?             8@        ������������������������       �                     @        �       �                    �?؇���X�?             5@        ������������������������       �                     $@        �       �                    �?���!pc�?             &@        ������������������������       �                      @        �       �                    �?�����H�?             "@        ������������������������       �                     @        �       �                    �N@z�G�z�?             @        ������������������������       �                     @        �       �                    �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?l��[B��?              M@       �       �                    �?����X�?             <@        ������������������������       �                     *@        �       �                    �?��S���?
             .@       �       �                   @b@�n_Y�K�?	             *@       �       �                   q@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �                          �^@�q�q�?             >@        ������������������������       �                      @                                �`@�eP*L��?	             6@                                �?�θ�?             *@       ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     "@        �t�bh�h)h,K ��h.��R�(KMKK��hb�BP  ZZZZZZ�?�������?��i��P�?����+�?�m۶m��?%I�$I��?*�Y7�"�?�����?      �?        9��8��?9��8���?�?�?              �?�q�q�?�q�q�?      �?      �?      �?                      �?              �?^Cy�5�?(������?      �?        �q�q�?�q�q�?              �?�������?�������?�q�q�?r�q��?              �?�������?�������?      �?              �?      �?      �?                      �?              �?R���Q�?ףp=
��?x6�;��?��
br�?�������?�������?�?�������?�$I�$I�?۶m۶m�?              �?      �?                      �?�%~F��?s��\;�?t�E]t�?]t�E�?x6�;��?��
br�?r�q��?�q�q�?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?O#,�4��?a���{�?              �?��(\���?{�G�z�?n۶m۶�?�$I�$I�?      �?        �������?�������?              �?      �?        F]t�E�?]t�E]�?      �?        �q�q�?9��8���?              �?      �?              �?        �$I�$I�?�m۶m��?      �?                      �?�������?�������?      �?        �������?�������?              �?      �?        n۶m۶�?%I�$I��?              �?�������?""""""�?F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?      �?              �?      �?              �?        y�5���?Cy�5��?F]t�E�?]t�E�?      �?      �?      �?                      �?              �?      �?      �?      �?        �������?�������?              �?      �?      �?              �?      �?        �ߔ�Ⱥ?	d����?���L�?�u�)�Y�?;�;��?ى�؉��?      �?        �q�q�?r�q��?              �?      �?        UUUUUU�?UUUUUU�?�?<<<<<<�?      �?      �?�$I�$I�?۶m۶m�?              �?      �?      �?              �?      �?                      �?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?        ہ�v`��?�g��%�?      �?      �?333333�?�������?              �?      �?        ^Cy�5�?(������?              �?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?      �?      �?      �?              �?      �?                      �?              �?              �?EQEQ�?�뺮��?�����?�����?M�[��?��'�W2�?�F�tj�?䮟-V��?d!Y�B�?�Mozӛ�?;ڼOqɐ?.�u�y�?              �?�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?      �?                      �?              �?L�Ϻ��?}���g�?�?�?�?<<<<<<�?              �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        F]t�E�?/�袋.�?�������?�������?      �?      �?      �?                      �?              �?      �?        q�f,��?<JeN���?�x+�R�?�Cj��V�?{�G�z�?
ףp=
�?              �?�a�a�?��y��y�?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?�������?�?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�����?���M���?2g�s��?sƜ1g̹?��8��8�?�q�q�?��F}g��?W�+�ɥ?��{���?�B!��?�����?8��18�?      �?      �?              �?      �?        >����?|���?      �?        <<<<<<�?�?UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?      �?        x����?����?|?_�_��?�A�A�?      �?        �������?�?      �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?      �?                      �?ffffff�?333333�?      �?      �?      �?                      �?      �?              �?      �?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        �������?ffffff�?      �?      �?�������?�������?              �?      �?                      �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?        F]t�E�?t�E]t�?              �?�q�q�?�q�q�?      �?        �������?�������?      �?              �?      �?              �?      �?        ���=��?GX�i���?�m۶m��?�$I�$I�?      �?        �������?�?ى�؉��?;�;��?t�E]t�?F]t�E�?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?              �?]t�E�?t�E]t�?ى�؉��?�؉�؉�?      �?                      �?              �?�t�bubhhubehhub.