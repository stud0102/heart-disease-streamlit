���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.3�ub�n_estimators�Kd�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhN�verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��Sex��ChestPainType��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��ExerciseAngina��Oldpeak��ST_Slope�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJV>rChG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h2�f8�����R�(KhONNNJ����J����K t�b�C              �?�t�bhSh&�scalar���hNC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hK�
node_count�K��nodes�h(h+K ��h-��R�(KK���h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(hh2�i8�����R�(KhONNNJ����J����K t�bK ��h�h�K��h�h�K��h�h_K��h�h_K ��h�h�K(��h�h_K0��uK8KKt�b�BX7         �                    �?��J�0�?=           ��@       u                    �?J3�xH��?9            �@       6       	          ����?�恾���?�            �v@                           �L@�Jhu4��?Y            @b@              	             ����*��?=            �X@������������������������       �                      @              
             �?�U�!��?<            @X@                          �n@�T|n�q�?            �E@	              	          833�?      �?             <@
                          �`@���}<S�?             7@������������������������       �                     1@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �        	             .@                          �b@�<ݚ�?"             K@                           @F@���B���?!             J@              	             �?�q�q�?             8@                           �?���N8�?             5@������������������������       �                     @������������������������       �        	             0@������������������������       �                     @                           �?@4և���?             <@������������������������       �                     6@                           T@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @       -                    �?��|�5��?            �G@       $                    _@      �?             @@        !                    �?���Q��?             @������������������������       �                     �?"       #       
             �?      �?             @������������������������       �                      @������������������������       �                      @%       (                    �?�>����?             ;@&       '                   f@      �?              @������������������������       �                     @������������������������       �                     �?)       *       	             �?�}�+r��?             3@������������������������       �                     0@+       ,       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @.       /                    �?��S���?	             .@������������������������       �                     @0       5                   p@���!pc�?             &@1       4                   @U@�����H�?             "@2       3       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @7       J                   `_@b<g���?            `k@8       E                    �?�>����?D             [@9       >                    �?(�5�f��?2            �S@:       =                    �M@"pc�
�?             &@;       <                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @?       D                    @I@ ��ʻ��?,             Q@@       C                    �? �q�q�?             8@A       B                   @[@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     5@������������������������       �                     F@F       I                    `@д>��C�?             =@G       H       
             �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     5@K       Z                    �?"��$�?;            �[@L       S                   �l@"pc�
�?             F@M       N       	             @��
ц��?             *@������������������������       �                     @O       P                     K@      �?              @������������������������       �                     @Q       R                     P@      �?             @������������������������       �                     �?������������������������       �                     @T       Y       	          ����?�g�y��?             ?@U       X                    �?�C��2(�?             &@V       W                    �N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        	             4@[       n                   0n@�iޤ��?&            �P@\       m       
             �?Hث3���?            �C@]       `                    �F@և���X�?            �A@^       _                    `@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@a       l                   �a@���|���?             6@b       k                    �?�z�G��?             4@c       f                   p`@ҳ�wY;�?
             1@d       e                   pj@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?g       h                    l@r�q��?             @������������������������       �                     @i       j                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @o       t                   �`@h�����?             <@p       s       	             �?z�G�z�?             @q       r                    �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     7@v       }                   x@BӀN��?a            �b@w       |                    �I@@ݚ)�?]             b@x       y       
             �?�Ra����?             F@������������������������       �                     ?@z       {                    b@�n_Y�K�?             *@������������������������       �                     @������������������������       �                      @������������������������       �        F             Y@~              	          ����?և���X�?             @������������������������       �                      @�       �                     L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   `@�iޤ��?            y@�       �                    �?j����?7            �T@�       �                    @JJ����?             �G@�       �                   �c@�Q����?             D@�       �                    �?z�G�z�?             4@�       �                    @K@�q�q�?             (@������������������������       �                     @�       �       	             �z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @L@R���Q�?             4@������������������������       �        	             "@�       �                    @P@���!pc�?             &@�       �                   �V@���Q��?             @������������������������       �                     �?�       �                   p@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �       	          033�?r�q��?             B@�       �       
             �?�����?             3@�       �                   �`@�r����?             .@�       �                   �[@�q�q�?             @������������������������       �                     @�       �                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     @������������������������       �        
             1@�       �       
             �?�f`��?�            �s@�       �                   �o@�A�|O��?G            @[@�       �                   ``@\I�~�?/            @S@�       �                   �e@�D��?            �H@�       �                    T@      �?             @@������������������������       �                     �?�       �                   `_@��a�n`�?             ?@�       �                    �? ��WV�?             :@������������������������       �                     5@�       �       	          `ff�?z�G�z�?             @�       �                   m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    `@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          033@��.k���?             1@�       �                   �Q@�q�q�?             (@������������������������       �                     @�       �                    �?�����H�?             "@�       �                   �e@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   ph@��X��?             <@�       �                   @e@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?��.k���?             1@�       �                    `P@��S���?
             .@�       �                    �?�n_Y�K�?	             *@������������������������       �                     @�       �                    �?X�<ݚ�?             "@�       �                   �c@����X�?             @�       �                   `l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                   �e@     ��?             @@�       �                    @K@¦	^_�?             ?@�       �                   �a@��S���?             .@������������������������       �                     @�       �       	             @�z�G��?             $@�       �                   `]@      �?              @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   Pr@      �?             0@������������������������       �        	             *@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    I@��
�j�?�            @j@�       �                   �`@      �?             @������������������������       �                      @�       �                    �?      �?             @�       �                    �F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   0h@`'�J�?�            �i@�       �                   �s@P����֨?�             i@�       �                    @L@ h'M#�?v            �f@������������������������       �        c            @c@�       �                    �? 	��p�?             =@�       �                   �l@z�G�z�?             $@������������������������       �                     @�       �                   �a@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     3@�       �                    @L@r�q��?
             2@������������������������       �                     *@�       �       	          ����?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�t�b�values�h(h+K ��h-��R�(KK�KK��h_�B�        x@     ��@      Z@     �y@      X@     �p@      N@     �U@     �H@      I@               @     �H@      H@      @      B@      @      5@       @      5@              1@       @      @       @                      @      @                      .@      E@      (@      E@      $@      0@       @      0@      @              @      0@                      @      :@       @      6@              @       @               @      @                       @      &@      B@      @      <@       @      @              �?       @       @               @       @               @      9@      �?      @              @      �?              �?      2@              0@      �?       @      �?                       @      @       @      @              @       @      �?       @      �?       @               @      �?                      @       @              B@     �f@       @      Y@      @      S@       @      "@       @       @       @                       @              @      �?     �P@      �?      7@      �?       @               @      �?                      5@              F@      @      8@      @      @      @                      @              5@      <@     �T@       @      B@      @      @              @      @      �?      @              @      �?              �?      @              �?      >@      �?      $@      �?      @              @      �?                      @              4@      4@     �G@      3@      4@      .@      4@      �?      (@      �?                      (@      ,@       @      ,@      @      &@      @      $@      �?      $@                      �?      �?      @              @      �?      �?              �?      �?              @                       @      @              �?      ;@      �?      @      �?       @      �?                       @               @              7@       @     �a@      @     `a@      @     �C@              ?@      @       @      @                       @              Y@      @      @       @              �?      @              @      �?             �q@      ^@      <@     �K@      6@      9@      5@      3@      @      0@      @       @              @      @      �?              �?      @                       @      1@      @      "@               @      @       @      @      �?              �?      @      �?                      @      @              �?      @      �?                      @      @      >@      @      *@       @      *@       @      @              @       @      �?              �?       @                      "@      @                      1@     �o@     @P@     �K@      K@     �F@      @@      B@      *@      <@      @              �?      <@      @      9@      �?      5@              @      �?       @      �?       @                      �?       @              @       @       @              �?       @              �?      �?      �?              �?      �?               @      "@       @      @              @       @      �?       @      �?              �?       @              @                      @      "@      3@      �?      $@              $@      �?               @      "@       @      @       @      @      @              @      @       @      @       @      �?       @                      �?              @       @                       @               @      $@      6@      "@      6@      @       @              @      @      @      @      �?       @      �?              �?       @              @                       @       @      ,@              *@       @      �?       @                      �?      �?             �h@      &@      @      @       @              �?      @      �?      �?      �?                      �?               @     �h@       @     �h@      @     �f@       @     @c@              ;@       @       @       @      @              @       @      @                       @      3@              .@      @      *@               @      @              @       @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJͥ�BhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK텔h~�B�3         �       
             �?<qn�h��?S           ��@                           �?j�q����?J           @@                          �c@�������?+             N@                          0c@x�K��?$            �I@                          �r@�[�IJ�?             �G@                          c@)O���?             B@                           �?J�8���?             =@       	                    �?l��
I��?             ;@������������������������       �        	             &@
                           �?      �?             0@                          �b@և���X�?             ,@                          �j@���Q��?	             $@������������������������       �                     @                          @b@և���X�?             @                           �?���Q��?             @              	          433�?      �?             @������������������������       �                     �?                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @                            K@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     @������������������������       �                     "@        �                    f@L��n��?           �{@!       0       	          ����?č�@��?           �z@"       /                    �L@h㱪��?E            �[@#       $                    �?�L#���?+            �P@������������������������       �                     I@%       &                    �?������?             1@������������������������       �                      @'       .                    �?�r����?
             .@(       )                   `]@z�G�z�?             $@������������������������       �                     @*       +                    �?���Q��?             @������������������������       �                     �?,       -                   `X@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                    �E@1       ^                    �?؇���X�?�            �s@2       =       
             �?N�zv�?>             V@3       4                    @I@��S���?
             .@������������������������       �                     @5       6                   �]@�q�q�?             (@������������������������       �                      @7       <       	          033@z�G�z�?             $@8       ;                   �`@�����H�?             "@9       :       	             @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?>       Q                   a@x�� ���?4            @R@?       @                   �_@��Q��?             D@������������������������       �        	             &@A       P                    �?l��[B��?             =@B       G                    �I@���|���?             6@C       D                    �?z�G�z�?             @������������������������       �                      @E       F                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @H       I                   Pl@������?             1@������������������������       �                     @J       K       	          `ff�?���|���?             &@������������������������       �                     @L       O                   Pb@z�G�z�?             @M       N                   m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @R       W                     Q@�C��2(�?            �@@S       T                    @h�����?             <@������������������������       �                     8@U       V                   �c@      �?             @������������������������       �                     �?������������������������       �                     @X       Y                    �?���Q��?             @������������������������       �                      @Z       ]                    �Q@�q�q�?             @[       \                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?_       ~                    �?0�N�]��?�            `l@`       i                   �[@�e�N�c�?{            �g@a       h                    �?���|���?
             6@b       c                   �W@�<ݚ�?	             2@������������������������       �                      @d       e       	          `ff�?      �?             0@������������������������       �                     $@f       g                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @j       s                   Xp@x�{�;��?q             e@k       r                   �c@�r�MȢ?G            �Z@l       q       	          ����?@䯦s#�?F            �Z@m       n                   �i@ �q�q�?             8@������������������������       �                     0@o       p                   �j@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �        5            �T@������������������������       �                     �?t       }                    �R@`Jj��?*             O@u       z                   0c@�.ߴ#�?)            �N@v       w                    �O@0�)AU��?&            �L@������������������������       �                     H@x       y                   ``@�����H�?             "@������������������������       �                     �?������������������������       �                      @{       |                     M@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?       �                    Y@r�q��?             B@������������������������       �                      @�       �                    @F@�t����?             A@������������������������       �                     �?�       �       	          ����?�C��2(�?            �@@�       �                   �l@����X�?             @������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @ ��WV�?             :@������������������������       �                     6@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @K@z�G�z�?	             .@�       �                   �`@$�q-�?             *@������������������������       �                     $@�       �                   @b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?VX����?	            z@�       �                   @E@��X�ە�?�            v@�       �                    �?J�8���?             =@�       �                    �?�z�G��?             4@�       �                   pb@��S�ۿ?
             .@������������������������       �        	             ,@������������������������       �                     �?������������������������       �                     @�       �                    ^@X�<ݚ�?             "@�       �       	             ��q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �? V䤾��?�            @t@�       �                   �a@�z�G��?-            �Q@������������������������       �                     9@�       �                    �?��S���?            �F@�       �                    �K@"pc�
�?             &@�       �                    �G@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �m@ҳ�wY;�?             A@�       �       	          033�?�q�����?             9@�       �                    b@�eP*L��?             6@�       �       	          ����?�q�q�?	             .@������������������������       �                     $@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                    @L@X�GP>��?�            �o@�       �                    �?�K��h�?~            �h@�       �                   �`@H%u��?             9@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @e@���7�?             6@������������������������       �                     5@������������������������       �                     �?������������������������       �        p            �e@�       �                    �?z�G�z�?"            �K@�       �                    �M@`2U0*��?             9@�       �                   �a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             5@�       �                   �^@�q�q�?             >@������������������������       �                      @�       �                   ps@X�Cc�?             <@�       �                    �? �o_��?             9@�       �                    d@      �?             0@�       �                    p@r�q��?
             (@������������������������       �                     @�       �                     M@���Q��?             @������������������������       �                     �?�       �                    @N@      �?             @�       �                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �p@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?^��>�b�?(            @P@������������������������       �                     &@�       �                    �?J��D��?#             K@�       �       	          ����?fP*L��?             F@�       �                    �?X�Cc�?
             ,@�       �                    p@      �?              @������������������������       �                     @�       �                   pq@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �a@      �?             @������������������������       �                     @������������������������       �                     @�       �                    @M@��S�ۿ?             >@������������������������       �                     &@�       �                    c@�KM�]�?             3@�       �       	          033�?�X�<ݺ?             2@������������������������       �        
             .@�       �                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       z@     P@     �V@     �y@      =@      ?@      4@      ?@      4@      ;@      3@      1@      3@      $@      3@       @      &@               @       @       @      @      @      @              @      @      @       @      @      �?      @              �?      �?       @               @      �?              �?               @              @                       @               @              @      �?      $@              $@      �?                      @      "@             �N@     �w@     �H@     �w@      @     �Z@      @     �O@              I@      @      *@       @               @      *@       @       @              @       @      @              �?       @       @       @                       @              @             �E@     �F@     �p@      9@     �O@       @      @              @       @      @               @       @       @       @      �?      @      �?      @                      �?      @                      �?      1@      L@      ,@      :@              &@      ,@      .@      ,@       @      �?      @               @      �?       @      �?                       @      *@      @      @              @      @      @              �?      @      �?      �?      �?                      �?              @              @      @      >@      �?      ;@              8@      �?      @      �?                      @       @      @               @       @      �?      �?      �?              �?      �?              �?              4@     �i@      ,@      f@       @      ,@      @      ,@       @               @      ,@              $@       @      @       @                      @      @              @     `d@       @     @Z@      �?     @Z@      �?      7@              0@      �?      @      �?                      @             �T@      �?              @      M@      @      M@      �?      L@              H@      �?       @      �?                       @       @       @               @       @              �?              @      >@       @              @      >@      �?              @      >@       @      @              @       @      �?              �?       @              �?      9@              6@      �?      @      �?                      @      (@      @      (@      �?      $@               @      �?              �?       @                       @     pt@     �V@     �r@      K@      $@      3@      @      ,@      �?      ,@              ,@      �?              @              @      @      @       @               @      @                      @     r@     �A@     �H@      5@      9@              8@      5@       @      "@       @      @              @       @                      @      6@      (@      *@      (@      $@      (@      $@      @      $@                      @              @      @              "@              n@      ,@     �h@      @      6@      @      �?       @      �?                       @      5@      �?      5@                      �?     �e@              F@      &@      8@      �?      @      �?              �?      @              5@              4@      $@       @              2@      $@      2@      @      $@      @      $@       @      @              @       @              �?      @      �?       @      �?              �?       @              �?                      @       @      �?       @                      �?              @      <@     �B@      &@              1@     �B@      @     �B@      @      "@       @      @              @       @      @       @                      @      @      @              @      @               @      <@              &@       @      1@      �?      1@              .@      �?       @      �?                       @      �?              $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJJ2:ihG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�Bx6         �       
             �?V�2���?5           ��@       k                   �b@l�,�Q�?C           H�@       2                    �?�3d`��?           �{@              	          ����?^��4m�?Z            �b@                          �X@ �h�7W�?!            �J@                          �W@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @	                           �F@`���i��?             F@
                           �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �C@       '                   �`@p�ݯ��?9            �W@       &                     Q@��S���?#             N@       %                   �b@|��?���?              K@              	          ����?�q�q�?             H@                           �M@z�G�z�?             4@                          �[@@4և���?             ,@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             &@              	             �?      �?             @������������������������       �                     @������������������������       �                     @                           @O@և���X�?             <@                          �a@z�G�z�?
             .@������������������������       �                     (@������������������������       �                     @                           �[@�	j*D�?             *@������������������������       �                      @!       $                    �?"pc�
�?             &@"       #       	          033�?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?������������������������       �                     @������������������������       �                     @(       +                   �]@z�G�z�?            �A@)       *                   `[@�eP*L��?             &@������������������������       �                     @������������������������       �                     @,       1                    �?�8��8��?             8@-       .       
             �?z�G�z�?             $@������������������������       �                     �?/       0                   �c@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@3       b                   �a@�F��O�?�            @r@4       S       	          ����?�*0��
�?�            `o@5       >                    �?��{H�?9            �U@6       7       	          ����?���|���?             &@������������������������       �                      @8       =                    �?�<ݚ�?             "@9       <                    �?      �?              @:       ;                   �e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �??       @       	          ����?@݈g>h�?1             S@������������������������       �                     :@A       F                   �Z@�:pΈ��?             I@B       C                   �_@����X�?             ,@������������������������       �                     "@D       E                    b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?G       H       	          `ff�?�8��8��?             B@������������������������       �                     $@I       L                    �L@ȵHPS!�?             :@J       K                   0a@�X�<ݺ?
             2@������������������������       �        	             1@������������������������       �                     �?M       N                   �]@      �?              @������������������������       �                     @O       P                    �?���Q��?             @������������������������       �                     �?Q       R                   8s@      �?             @������������������������       �                      @������������������������       �                      @T       Y                   �b@��Y��]�?f            �d@U       V                    �? 4^��?K            �]@������������������������       �        >            �X@W       X                    �?P���Q�?             4@������������������������       �                     �?������������������������       �                     3@Z       _                   �_@��S�ۿ?            �F@[       ^       
             �?�?�|�?            �B@\       ]                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     >@`       a                   `@      �?              @������������������������       �                      @������������������������       �                     @c       j                   �k@�p ��?            �D@d       i                    �J@      �?             (@e       h                   i@�q�q�?             "@f       g                     I@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     =@l       �                   �o@�5��?3            @T@m       n                   @J@�E��ӭ�?!             K@������������������������       �                      @o       z                   0d@      �?              J@p       q                    @C@؇���X�?             <@������������������������       �                     �?r       w       	             @�����H�?             ;@s       v                   �g@ �q�q�?             8@t       u                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@x       y                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @{       �       	          ����?      �?             8@|       }                   @_@      �?             0@������������������������       �                     $@~       �                   �`@�q�q�?             @       �                    f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                      @�       �                   g@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �e@�q�q�?             ;@�       �                   �`@��<b���?             7@������������������������       �                     (@�       �                    @�eP*L��?             &@�       �                    q@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�ၝ���?�            �x@�       �                    c@�MI8d�?�            �t@�       �                    �?F�����?            �F@�       �                   �b@�q�q�?             8@�       �                    _@��s����?             5@�       �                   @\@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?@4և���?             ,@������������������������       �                     &@�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     5@�       �                   �g@�5?,R�?�             r@�       �                    �?@2����?�            �q@�       �                    �M@`2U0*��?A             Y@������������������������       �        2            @R@�       �                   �r@PN��T'�?             ;@������������������������       �        	             .@�       �                   d@�q�q�?             (@������������������������       �                      @������������������������       �                     @�       �                   �h@��r
'��?l            @g@������������������������       �                     C@�       �       	          ����?$G$n��?X            �b@�       �                    ]@@���|N�?M             `@�       �                    �?     ��?             @@�       �                   �[@���Q��?             @�       �                   Pa@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   �b@�����H�?             ;@������������������������       �                     *@�       �                   @c@d}h���?             ,@������������������������       �                      @�       �                    �?�8��8��?             (@�       �                    �H@�C��2(�?             &@������������������������       �                      @�       �                    �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �t@��8�$>�?<            @X@�       �                    @N@��<b�ƥ?8             W@�       �                    �?���E�?4            �U@�       �                   0e@�}�+r��?
             3@������������������������       �                     .@�       �                    �H@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        *             Q@�       �                   pj@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   u@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    b@�\��N��?             3@�       �                   ``@r�q��?             (@�       �                   xp@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �]@      �?)             P@�       �                     K@����X�?             ,@������������������������       �                     @������������������������       �                     $@�       �                    d@� �	��?!             I@�       �                    �?�q�q�?             B@������������������������       �                     @�       �                    �?     ��?             @@�       �                   �`@      �?             <@�       �                    �?���Q��?             .@�       �                    n@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   0a@X�<ݚ�?             "@�       �                   �_@�q�q�?             @�       �                    �?z�G�z�?             @�       �                   �l@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �H@$�q-�?             *@������������������������       �                      @�       �                   `j@z�G�z�?             @������������������������       �                     @�       �                    @J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   Pe@@4և���?             ,@������������������������       �                      @�       �                    �G@r�q��?             @������������������������       �                      @�       �                   pf@      �?             @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       Pz@     @     �[@     �y@      O@     �w@      C@     �[@      @      I@       @      @              @       @              �?     �E@      �?      @      �?                      @             �C@     �A@      N@      <@      @@      <@      :@      <@      4@      0@      @      *@      �?       @      �?       @                      �?      &@              @      @      @                      @      (@      0@      @      (@              (@      @              "@      @               @      "@       @      "@      �?              �?      "@                      �?              @              @      @      <@      @      @              @      @               @      6@       @       @      �?              �?       @               @      �?                      ,@      8@     �p@      2@      m@      ,@     @R@      @      @               @      @       @      @      �?       @      �?       @                      �?      @                      �?      @     @Q@              :@      @     �E@      @      $@              "@      @      �?      @                      �?      @     �@@              $@      @      7@      �?      1@              1@      �?               @      @              @       @      @              �?       @       @               @       @              @      d@      �?     �]@             �X@      �?      3@      �?                      3@      @      E@      �?      B@      �?      @              @      �?                      >@       @      @       @                      @      @     �A@      @      @      @      @       @      @              @       @              @                      @              =@      H@     �@@     �C@      .@               @     �C@      *@      8@      @              �?      8@      @      7@      �?      �?      �?      �?                      �?      6@              �?       @      �?                       @      .@      "@      (@      @      $@               @      @      �?      @              @      �?              �?              @      @       @              �?      @              @      �?              "@      2@      @      2@              (@      @      @      @      @              @      @                      @      @             ps@     �U@     pq@      K@      1@      <@      1@      @      1@      @      @      @      @                      @      *@      �?      &@               @      �?              �?       @                      @              5@     `p@      :@     `p@      8@      X@      @     @R@              7@      @      .@               @      @       @                      @     �d@      4@      C@              `@      4@     �]@      $@      :@      @       @      @       @       @       @                       @              �?      8@      @      *@              &@      @               @      &@      �?      $@      �?       @               @      �?              �?       @              �?             @W@      @     �V@       @     �U@      �?      2@      �?      .@              @      �?              �?      @              Q@              @      �?              �?      @              @       @               @      @              "@      $@       @      $@       @      @              @       @                      @      @                       @      @@      @@      @      $@      @                      $@      <@      6@      .@      5@      @              &@      5@      @      5@      @      "@      �?      @      �?                      @      @      @       @      @      �?      @      �?      @              @      �?                      �?      �?              @              �?      (@               @      �?      @              @      �?      �?      �?                      �?      @              *@      �?       @              @      �?       @              @      �?              �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJH��0hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM#hwh(h+K ��h-��R�(KM#��h~�B�?         �                    �?>���i��?M           ��@       )                    �?0����;�?H           �@                          �R@:2vz�M�?-            �N@������������������������       �                      @                           �?�F�j��?(            �J@              	          `ff@��+7��?             7@                          �b@��s����?             5@       	       	          ����?@4և���?
             ,@������������������������       �                     "@
                          �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                           �I@և���X�?             @������������������������       �                      @                          p@���Q��?             @������������������������       �                     �?                          �b@      �?             @                          �v@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                          �q@�z�G��?             >@                          @n@��S�ۿ?             .@������������������������       �                     @                            I@      �?              @                          �n@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       "                    @L@��S���?             .@        !                   �_@r�q��?             @������������������������       �                     �?������������������������       �                     @#       (                    �?�<ݚ�?             "@$       %       	          ����?      �?              @������������������������       �                     @&       '                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?*       q       	          033�?B�&��*�?           �{@+       4                   @E@>��"��?n            �e@,       3                    @N@�:�]��?             �I@-       .       
             �?��-�=��?            �C@������������������������       �                     ;@/       2                    �?�q�q�?             (@0       1                   @_@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     (@5       X                   ``@N1���?N            �^@6       Q                    �?^�JB=�?1            @T@7       P                    �?�m����?$            �M@8       E                   �b@���H.�?              I@9       D                    @K@�>4և��?             <@:       ?                   ``@X�Cc�?             ,@;       <                   �Z@�q�q�?             @������������������������       �                     �?=       >                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?@       C                   �l@      �?              @A       B                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@F       G                    �B@���!pc�?             6@������������������������       �                      @H       O                   �p@z�G�z�?             4@I       N                   �n@���Q��?             $@J       K                   @^@      �?              @������������������������       �                     @L       M                   �j@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     $@������������������������       �                     "@R       S                    @N@�C��2(�?             6@������������������������       �        	             0@T       U                    �?�q�q�?             @������������������������       �                     @V       W                    �P@�q�q�?             @������������������������       �                      @������������������������       �                     �?Y       f                   �a@hP�vCu�?            �D@Z       a       
             �?�θ�?             :@[       ^                   0a@      �?              @\       ]                    q@z�G�z�?             @������������������������       �                     �?������������������������       �                     @_       `                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @b       e                   �f@�X�<ݺ?             2@c       d                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             0@g       p       	             �?�q�q�?             .@h       o                     M@�n_Y�K�?             *@i       n                   �e@����X�?             @j       k                    b@r�q��?             @������������������������       �                      @l       m       
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @r       s                   �U@���x���?�            �p@������������������������       �                     �?t       �                   Pf@�\�)G�?�            �p@u       �                   pv@�qM�R��?�            �p@v       �                   pb@$�q-�?�            @p@w       �                    �?P���Q�?�             i@x       �                    �O@`-�I�w�?a             c@y       �       	             �?6uH���?O             _@z       �                    �?�t����?             A@{       |                   ``@$�q-�?             :@������������������������       �                     ,@}       ~                   �m@r�q��?
             (@������������������������       �                     @       �                    @K@�q�q�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �X@      �?              @������������������������       �                     �?�       �                    ^@؇���X�?             @�       �                   �Y@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �Z@��S�ۿ?8            �V@�       �                   �X@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �T@Pq�����?6            @U@�       �                    �L@����X�?             @������������������������       �                     @������������������������       �                      @�       �                   �\@ ���J��?2            �S@�       �       	             �?ףp=
�?             $@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    @M@ ��ʻ��?,             Q@������������������������       �                     G@�       �                    �M@���7�?             6@�       �       	          `ff�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     3@������������������������       �                     <@������������������������       �        $             H@�       �                    �?r�q��?"             N@�       �                     P@X�Cc�?             ,@������������������������       �                     @�       �       
             �?����X�?             @������������������������       �                      @������������������������       �                     @�       �                   �e@�q��/��?             G@�       �                    c@���Q��?             $@�       �                   �Z@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �r@������?             B@������������������������       �                     ;@�       �                    �R@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                   �|@      �?              @�       �                   `a@z�G�z�?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       
             �?��ۉ���?           �y@�       �                   p`@��u����?]             c@�       �       	          ����?��q7L��?0            �T@�       �       
             �?؇���X�?
             ,@������������������������       �                     �?�       �                    �J@$�q-�?	             *@�       �                    �F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@�       �                    �?��z4���?&            @Q@�       �                   @[@����X�?             <@������������������������       �                      @�       �                   `m@�θ�?             :@�       �                   `b@��
ц��?             *@�       �                     R@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �K@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@�       �                    �?�>$�*��?            �D@�       �                   @c@���Q��?             @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   `k@�q�q�?             B@�       �       	             @      �?	             0@������������������������       �                     *@�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    f@��Q��?             4@�       �                   �c@��S���?	             .@�       �       	          `ff�?�q�q�?             (@�       �                    @z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?4�2%ޑ�?-            �Q@�       �       	          ����?���Q��?
             .@�       �                   @a@      �?              @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    `@X�;�^o�?#            �K@������������������������       �                     :@�       �       	          833�?>���Rp�?             =@�       �                    �?���Q��?             @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �a@r�q��?             8@������������������������       �                     *@�       �                    �M@���|���?             &@������������������������       �                     @�       �       	          hff�?      �?              @������������������������       �                      @�       �                    `P@�q�q�?             @������������������������       �                     @������������������������       �                      @�                           X@P�� �?�            @p@������������������������       �                      @      "      	             @x�]AgȽ?�             p@            	            �?�nkK�?�            �o@                        �s@ f^8���?�            �i@      	                  @[@�q�q�?{             h@                         �?@4և���?
             ,@������������������������       �                     &@                        `^@�q�q�?             @������������������������       �                      @������������������������       �                     �?
                        �c@@~��?q            @f@������������������������       �        f            �c@                        �d@���N8�?             5@                        `R@@4և���?             ,@������������������������       �                     �?������������������������       �                     *@������������������������       �                     @                        �`@����X�?	             ,@������������������������       �                     "@                        �a@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                         �?�*/�8V�?             �G@                         @L@@4և���?             E@������������������������       �                     ?@                        @b@���!pc�?             &@                        �`@      �?             @������������������������       �                      @������������������������       �                      @                        �k@؇���X�?             @������������������������       �                     �?������������������������       �                     @       !                  �b@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�t�b��0     h�h(h+K ��h-��R�(KM#KK��h_�B0       �y@     �@     @\@     �x@      :@     �A@               @      :@      ;@      1@      @      1@      @      *@      �?      "@              @      �?      @                      �?      @      @       @               @      @      �?              �?      @      �?      �?              �?      �?                       @               @      "@      5@      �?      ,@              @      �?      @      �?      �?      �?                      �?              @       @      @      �?      @      �?                      @      @       @      @      �?      @               @      �?              �?       @                      �?     �U@     Pv@      N@     @\@      @     �G@      @     �A@              ;@      @       @      @      @              @      @                      @              (@      L@     �P@      ?@      I@      =@      >@      =@      5@      7@      @      "@      @       @      @      �?              �?      @              @      �?              @      �?       @      �?       @                      �?      @              ,@              @      0@       @              @      0@      @      @       @      @              @       @      �?              �?       @               @                      $@              "@       @      4@              0@       @      @              @       @      �?       @                      �?      9@      0@      4@      @      @      @      �?      @      �?                      @       @      �?              �?       @              1@      �?      �?      �?      �?                      �?      0@              @      $@      @       @      @       @      @      �?       @              @      �?              �?      @                      �?              @               @      ;@     �n@      �?              :@     �n@      8@     �n@      4@      n@      $@     �g@      $@     �a@      $@     �\@      @      >@       @      8@              ,@       @      $@              @       @      @       @      �?              �?       @                      @       @      @      �?              �?      @      �?       @               @      �?                      @      @      U@       @      @              @       @              @     @T@       @      @              @       @               @      S@      �?      "@      �?       @               @      �?                      @      �?     �P@              G@      �?      5@      �?       @               @      �?                      3@              <@              H@      $@      I@      @      "@              @      @       @               @      @              @     �D@      @      @      @      �?              �?      @                      @      �?     �A@              ;@      �?       @               @      �?              @      @      @      �?       @               @      �?       @                      �?              @       @             �r@     �\@      L@     @X@      D@     �E@       @      (@      �?              �?      (@      �?       @               @      �?                      $@      C@      ?@      4@       @               @      4@      @      @      @      @      �?      @                      �?      �?      @      �?                      @      *@              2@      7@      @       @      �?       @               @      �?               @              .@      5@       @      ,@              *@       @      �?       @                      �?      *@      @       @      @       @      @       @       @       @                       @               @              @      @              0@      K@      "@      @       @      @       @      �?              �?       @                      @      @              @      H@              :@      @      6@      @       @       @              �?       @      �?                       @      @      4@              *@      @      @              @      @      @               @      @       @      @                       @     @n@      2@               @     @n@      0@     @n@      &@      i@      @     �g@       @      *@      �?      &@               @      �?       @                      �?      f@      �?     �c@              4@      �?      *@      �?              �?      *@              @              $@      @      "@              �?      @              @      �?              E@      @     �C@      @      ?@               @      @       @       @               @       @              @      �?              �?      @              @       @               @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ$��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B88         �                    �?&�L�m��?L           ��@       ?                    �?,���0�?3           �}@       4                    �?��k4C��?            �h@              
             �?JJ����?Y            �a@       
                    �?����>4�?'             L@       	                   �b@      �?
             ,@                          �a@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @                          �e@�����?             E@                           �?��p\�?            �D@                          �^@��?^�k�?            �A@                           @H@�C��2(�?             &@������������������������       �                     @                          �p@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     8@              	             �?�q�q�?             @������������������������       �                      @                           `@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?                           �?f��>���?2            @U@                           s@ףp=
�?             4@������������������������       �        
             2@������������������������       �                      @       %                    �?R=6�z�?&            @P@       $                   �a@�q�q�?             (@        #                   �\@z�G�z�?             $@!       "                    `@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @&       1       	            �? {��e�?             �J@'       .                   �b@ >�֕�?            �A@(       -                    ]@Pa�	�?            �@@)       *                   �b@r�q��?             @������������������������       �                     @+       ,                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ;@/       0                    �?      �?              @������������������������       �                     �?������������������������       �                     �?2       3                   P`@      �?             2@������������������������       �                     "@������������������������       �                     "@5       6       
             �? 	��p�?&             M@������������������������       �                     F@7       >       	          ����?����X�?	             ,@8       9       	          ,33ӿ      �?              @������������������������       �                     @:       ;                    �?z�G�z�?             @������������������������       �                     @<       =                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @@       O       	          hff�?�ܸb���?�            @q@A       B                   �i@�q�q�?             H@������������������������       �        	             1@C       N                   @e@�4�����?             ?@D       M                   `a@      �?             <@E       L                   �d@p�ݯ��?             3@F       I                   8p@      �?
             0@G       H                   �`@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?J       K       	          ����?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     "@������������������������       �                     @P       �                    �?`� x��?�            �l@Q       R                   �U@�T_�/��?p            `d@������������������������       �                      @S       t       	          ����?������?o             d@T       i       	          033�?v���a�?2            @R@U       h                   ``@lGts��?&            �K@V       Y                    �H@�MI8d�?            �B@W       X                   `o@�q�q�?             @������������������������       �                      @������������������������       �                     �?Z       g                   @e@�t����?             A@[       ^       	          ����?�C��2(�?            �@@\       ]                    Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?_       `                    �?��S�ۿ?             >@������������������������       �                     �?a       f                   �X@XB���?             =@b       e                   l@r�q��?             @c       d                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     7@������������������������       �                     �?������������������������       �                     2@j       q                    �?�E��ӭ�?             2@k       l                   @]@d}h���?	             ,@������������������������       �                     @m       n                     I@      �?              @������������������������       �                     @o       p                   �`@      �?             @������������������������       �                     @������������������������       �                     �?r       s                   @[@      �?             @������������������������       �                      @������������������������       �                      @u       �                   `q@���7�?=             V@v       }                    �?,�+�C�?(            �K@w       |                   q@���N8�?             E@x       y       
             �?��Y��]�?            �D@������������������������       �                    �C@z       {                   `W@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?~                            K@8�Z$���?	             *@������������������������       �                      @������������������������       �                     &@������������������������       �                    �@@������������������������       �        *            @P@�       �       
             �?����W��?           �{@�       �                   �b@"�!���?n            �d@�       �                    �?r�z-��?H            �Z@�       �                   @_@��>4և�?             <@�       �       	          ���ɿףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �?X�<ݚ�?             2@�       �                   �k@�q�q�?             (@�       �       	          833�?      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �n@      �?              @������������������������       �                     @�       �                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �R@����?7            �S@�       �                   �e@N��c��?6            @S@�       �                    �?�>����?             ;@�       �       
             �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�nkK�?             7@�       �                    @L@�����H�?             "@�       �       	             �r�q��?             @������������������������       �                     @�       �                    @K@�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        
             ,@�       �                    �?`�Q��?"             I@�       �                   @Z@hP�vCu�?            �D@������������������������       �                      @�       �                    �?�99lMt�?            �C@�       �       	          @33�?     ��?             @@�       �                   �`@ףp=
�?             $@�       �                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �b@���|���?             6@�       �                    @F@��S���?             .@������������������������       �                     @�       �                    �?�q�q�?
             (@�       �                    @�q�q�?             @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   @q@؇���X�?             @�       �                   �o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   pb@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     �?�       �                    �F@��6}��?&            �N@�       �                    @P���Q�?             4@������������������������       �        
             3@������������������������       �                     �?�       �       	          ����?��]�T��?            �D@�       �                    @      �?              @�       �                   �p@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   Pc@���!pc�?            �@@������������������������       �                      @�       �                   �c@��H�}�?             9@������������������������       �                     @�       �                   �l@���N8�?             5@������������������������       �                     "@�       �                   Pr@�q�q�?	             (@�       �       	          ���@      �?              @�       �                    �?����X�?             @������������������������       �                     �?�       �       	          ����?r�q��?             @�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �O@Xe�&��?�            @q@�       �                   Pa@j���� �?
             1@�       �                   `X@����X�?             ,@������������������������       �                      @�       �       	          ����?r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     @�       �                   �p@ 8i%M�?�            0p@�       �                    �L@     ��?w             h@�       �                    @G@��ϩ}��?g            �d@������������������������       �        6             V@�       �                    �G@�e���@�?1            @S@�       �                    o@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        -            �Q@�       �                   `l@�>����?             ;@�       �                    @r�q��?             (@�       �                   �`@�C��2(�?             &@�       �                   @`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     .@�       �                    �?pH����?*            �P@������������������������       �                    �A@�                           �?     ��?             @@�       �                   c@\-��p�?             =@������������������������       �                     8@�       �                   `r@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�B       �{@     �}@     �Z@     w@     �S@      ^@     �R@     �P@      &@     �F@      @      @      @      @      @                      @              @      @      C@      @      C@      �?      A@      �?      $@              @      �?      @              @      �?                      8@       @      @               @       @       @       @                       @      �?              P@      5@      2@       @      2@                       @      G@      3@      @       @       @       @       @      @       @                      @              @       @              E@      &@     �@@       @      @@      �?      @      �?      @              �?      �?      �?                      �?      ;@              �?      �?              �?      �?              "@      "@              "@      "@              @      K@              F@      @      $@      @      @              @      @      �?      @              �?      �?              �?      �?                      @      ;@      o@      $@      C@              1@      $@      5@      @      5@      @      (@      @      (@      �?      $@              $@      �?              @       @               @      @              @                      "@      @              1@     `j@      1@     @b@       @              .@     @b@      &@      O@      @     �H@      @      ?@       @      �?       @                      �?      @      >@      @      >@      �?       @               @      �?               @      <@      �?              �?      <@      �?      @      �?      �?      �?                      �?              @              7@      �?                      2@      @      *@      @      &@              @      @      @              @      @      �?      @                      �?       @       @       @                       @      @      U@      @     �I@       @      D@      �?      D@             �C@      �?      �?      �?                      �?      �?               @      &@       @                      &@             �@@             @P@     @u@     �Y@     @T@     �U@      B@     �Q@      1@      &@      "@      �?              �?      "@               @      $@       @      @      �?      @              @      �?              @      �?      @               @      �?              �?       @                      @      3@     �M@      2@     �M@       @      9@      �?      @      �?                      @      �?      6@      �?       @      �?      @              @      �?       @              �?      �?      �?      �?                      �?              @              ,@      0@      A@      0@      9@       @              ,@      9@      "@      7@      �?      "@      �?       @               @      �?                      @       @      ,@      @       @      @              @       @      @       @      �?       @               @      �?              @                      @      �?      @      �?      �?              �?      �?                      @      @       @               @      @                      "@      �?             �F@      0@      3@      �?      3@                      �?      :@      .@       @      @      �?      @              @      �?              �?              8@      "@       @              0@      "@              @      0@      @      "@              @      @      @      @       @      @      �?              �?      @      �?      �?      �?                      �?              @      �?              @             0p@      1@      $@      @      $@      @               @      $@       @      $@                       @              @      o@      $@     �g@      @     �d@      �?      V@              S@      �?      @      �?              �?      @             �Q@              9@       @      $@       @      $@      �?      @      �?      @                      �?      @                      �?      .@              N@      @     �A@              9@      @      9@      @      8@              �?      @              @      �?                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ(�*RhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�7         �                    �?TU�`��?Q           ��@       q                    �?�+d����?�           ��@       8                    �?pa���i�?�            �u@                           �?\��_��?[            �a@       
                    b@�θ�?            �C@                          �s@�g�y��?             ?@������������������������       �                     ;@       	                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @       -                   �`@������?B            �Y@                          @E@:-�.A�?.            �P@              
             �?      �?	             0@������������������������       �                     @                           �?�����H�?             "@                           �G@z�G�z�?             @������������������������       �                      @              	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @       *                    �?ҳ�wY;�?%            �I@              
             �?�X����?             F@              	          ����?H%u��?             9@������������������������       �                     1@                           �F@      �?              @������������������������       �                      @                          `a@r�q��?             @������������������������       �                     @������������������������       �                     �?        #                    �?D�n�3�?             3@!       "                   �f@z�G�z�?             @������������������������       �                     @������������������������       �                     �?$       )       	          hff�?����X�?             ,@%       &                    �I@r�q��?
             (@������������������������       �                     @'       (                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @+       ,       
             �?և���X�?             @������������������������       �                     @������������������������       �                     @.       3       
             �?      �?             B@/       2                    �L@���!pc�?             &@0       1       	          ����?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @4       5                    @N@`2U0*��?             9@������������������������       �                     7@6       7                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?9       p                   pf@,���i�?�            �i@:       ;                   �U@pH����?�             i@������������������������       �                     @<       o       	          `ff @�C��2(�?�            �h@=       N                    �?�q��/��?^            `b@>       M                    f@�E��ӭ�?             2@?       B                   �`@������?             1@@       A       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?C       L                   �a@؇���X�?
             ,@D       G       	             �?      �?              @E       F                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?H       I                    �I@r�q��?             @������������������������       �                     @J       K                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?O       T                    @J@�|K��2�?P             `@P       Q                   pb@h�����?             L@������������������������       �                    �E@R       S                     E@8�Z$���?             *@������������������������       �                      @������������������������       �                     &@U       n                   (q@v���a�?3            @R@V       k                   �b@����>4�?)             L@W       b       	          hff�?L紂P�?'            �I@X       Y                   `Y@�<ݚ�?             2@������������������������       �                     @Z       ]                   @\@����X�?
             ,@[       \                    k@���Q��?             @������������������������       �                      @������������������������       �                     @^       a                   �T@�����H�?             "@_       `                     P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @c       j                   �i@�C��2(�?            �@@d       e                   �\@r�q��?             2@������������������������       �                     �?f       i                    I@�t����?             1@g       h                   `_@"pc�
�?	             &@������������������������       �                     "@������������������������       �                      @������������������������       �                     @������������������������       �                     .@l       m       
             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             1@������������������������       �        "            �I@������������������������       �                     @r       �                    @L@>��C��?�            �u@s       �       
             �?���O1��?�             o@t       w                    �?     ��?+             P@u       v                    V@�����H�?             "@������������������������       �                     �?������������������������       �                      @x       �                    �K@N{�T6�?#            �K@y       �                    �E@�q�q�?!            �I@z       {                   pf@���!pc�?             &@������������������������       �                     �?|              	          033@z�G�z�?             $@}       ~                    @�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �q@R���Q�?             D@�       �                    @J@�z�G��?             >@�       �                   @m@z�G�z�?             4@�       �                    �?�t����?             1@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @^@@4և���?	             ,@�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                   e@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �K@      �?             $@������������������������       �                     �?�       �                    �?X�<ݚ�?             "@�       �       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     @�       �       	             �? S5W�?�             g@������������������������       �        t            �d@�       �                    �?�X�<ݺ?             2@�       �                   `^@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       �       
             �?���̅��?=            �W@�       �                   Pg@(���@��?            �G@�       �                    �P@�r����?             .@������������������������       �                     "@�       �       
             �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �O@     ��?             @@�       �                    Y@�GN�z�?             6@������������������������       �                     �?�       �                    \@��s����?             5@������������������������       �                      @�       �                    �N@�KM�]�?             3@�       �                    �?      �?
             0@�       �                    @M@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �P@z�G�z�?             $@������������������������       �                     @�       �                   pj@      �?             @������������������������       �                      @������������������������       �                      @�       �       	          ��� @      �?             H@�       �                    �L@��|�5��?            �G@������������������������       �                     @�       �                   �j@"pc�
�?             F@�       �                   �h@���Q��?
             .@�       �                    �?"pc�
�?	             &@������������������������       �                     @�       �                    `Q@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	          ����? 	��p�?             =@�       �                    �?�r����?	             .@�       �                   pb@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   ps@�8��8��?             (@������������������������       �                     $@�       �                   u@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             ,@������������������������       �                     �?�       �       	          ����?�G��6�?�            `l@�       �                   �O@�����?9            �V@������������������������       �                    �D@�       �                    �?z�):���?!             I@�       �       
             �?��s����?             5@������������������������       �        
             1@������������������������       �                     @�       �                   �W@V�a�� �?             =@������������������������       �                     �?�       �                   �d@�>4և��?             <@�       �       
             �?��<b���?             7@�       �                   `c@z�G�z�?             @������������������������       �                     @�       �                     P@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�X�<ݺ?             2@�       �                    �?z�G�z�?             @�       �                   o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     @�       �                    �?l��\��?R             a@�       �                    �?@��,B�?:            �V@�       �                   @Y@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        6            @U@�       �                   Pb@��Hg���?            �F@�       �                   pb@�IєX�?             A@������������������������       �                     ?@�       �                   `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @H@"pc�
�?	             &@�       �                     F@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	             @�����H�?             "@������������������������       �                     @�       �                    �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       @y@     �@     �v@     `t@     @Y@     �n@      S@     �P@      >@      "@      >@      �?      ;@              @      �?              �?      @                       @      G@     �L@      3@      H@      �?      .@              @      �?       @      �?      @               @      �?       @      �?                       @              @      2@     �@@      ,@      >@      @      6@              1@      @      @       @              �?      @              @      �?              &@       @      �?      @              @      �?              $@      @      $@       @      @              @       @               @      @                       @      @      @              @      @              ;@      "@      @       @      @       @               @      @                      @      8@      �?      7@              �?      �?      �?                      �?      9@     �f@      5@     �f@      @              2@     �f@      2@      `@      @      *@      @      *@       @      �?       @                      �?       @      (@       @      @      �?      �?              �?      �?              �?      @              @      �?      �?              �?      �?                      @      �?              *@      ]@       @      K@             �E@       @      &@       @                      &@      &@      O@      &@     �F@      @      F@      @      ,@              @      @      $@      @       @               @      @              �?       @      �?      �?      �?                      �?              @      @      >@      @      .@      �?               @      .@       @      "@              "@       @                      @              .@      @      �?      @                      �?              1@             �I@      @             �p@      T@     �j@      B@      =@     �A@       @      �?              �?       @              5@      A@      1@      A@       @      @              �?       @       @       @      �?       @                      �?              �?      "@      ?@      "@      5@      @      0@       @      .@      �?       @               @      �?              �?      *@      �?       @      �?                       @              &@       @      �?       @                      �?      @      @              �?      @      @      @       @               @      @              �?       @      �?                       @              $@      @              g@      �?     �d@              1@      �?      @      �?              �?      @              (@             �I@      F@      .@      @@       @      *@              "@       @      @              @       @              *@      3@      @      1@      �?              @      1@       @               @      1@      �?      .@      �?      @              @      �?                      &@      �?       @               @      �?               @       @      @               @       @       @                       @      B@      (@      B@      &@              @      B@       @      "@      @      "@       @      @               @       @       @                       @              @      ;@       @      *@       @       @      �?       @                      �?      &@      �?      $@              �?      �?              �?      �?              ,@                      �?     �C@     �g@      ;@      P@             �D@      ;@      7@      @      1@              1@      @              7@      @              �?      7@      @      2@      @      �?      @              @      �?      �?              �?      �?              1@      �?      @      �?       @      �?       @                      �?       @              *@              @              (@      _@      �?     �V@      �?      @      �?                      @             @U@      &@      A@       @      @@              ?@       @      �?       @                      �?      "@       @      �?      �?      �?                      �?       @      �?      @               @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���}hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM	hwh(h+K ��h-��R�(KM	��h~�B�9         �       
             �?T �����?N           ��@       w                   Pb@�㙢�c�?M           �@       J                    �?HX���?           �x@       	                   `[@�x`a��?�            s@              	          hff�?��'�`�?6            �T@              	          ����?P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �        (            �O@
       %                   �_@̹�"���?�            �k@                           \@r�q��?-            �P@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @       $                   `_@�?�P�a�?*             N@                          @^@��ϭ�*�?)             M@������������������������       �        
             .@                          �h@X�EQ]N�?            �E@������������������������       �                     5@              
             �?�GN�z�?             6@������������������������       �                     @       #       	             �?�E��ӭ�?             2@       "       	          ����?�eP*L��?             &@                           �?�q�q�?             "@������������������������       �                     �?       !       	          ����?      �?              @                            �?�q�q�?             @                          q@z�G�z�?             @������������������������       �                     @                           @D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @&       '                    �?��)�G��?d            �c@������������������������       �                     B@(       A                   `@�.�?�P�?O             ^@)       ,                    �?�r����?3            �R@*       +                   �_@      �?              @������������������������       �                     @������������������������       �                     @-       <                   `_@pH����?.            �P@.       1                   �[@����˵�?(            �M@/       0       	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @2       9                    �R@ 7���B�?#             K@3       8                    �? pƵHP�?!             J@4       5                   �p@r�q��?             @������������������������       �                     @6       7                   hs@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     G@:       ;       	             @      �?              @������������������������       �                     �?������������������������       �                     �?=       >                    �?      �?              @������������������������       �                     �??       @                    �F@և���X�?             @������������������������       �                     @������������������������       �                     @B       I                    �?����?�?            �F@C       D                    �?@4և���?             ,@������������������������       �                     @E       H                   �m@ףp=
�?             $@F       G                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     ?@K       f                   0`@      �??             V@L       c       	          `ff@     ��?-             P@M       b                    �R@�?�P�a�?+             N@N       a                    �?��ϭ�*�?*             M@O       ^                    `Q@,���i�?            �D@P       ]                   P`@�L���?            �B@Q       Z       	          `ff�?r�q��?             2@R       Y                   �_@@4և���?	             ,@S       X                    �?�����H�?             "@T       U                    �?�q�q�?             @������������������������       �                     �?V       W                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @[       \       	          033�?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     3@_       `                   �Z@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     1@������������������������       �                      @d       e                    �?      �?             @������������������������       �                     �?������������������������       �                     @g       r                   o@      �?             8@h       i                    �?ҳ�wY;�?             1@������������������������       �                     @j       q                    �?      �?	             (@k       p                     Q@�eP*L��?             &@l       m                   �j@X�<ݚ�?             "@������������������������       �                     @n       o                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?s       t                   �p@؇���X�?             @������������������������       �                     @u       v                   pq@      �?              @������������������������       �                     �?������������������������       �                     �?x       �                    �?�ݧ�N,�?G            @\@y       ~                    �G@8��8���?             H@z       }                    �?      �?             0@{       |                   @q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@       �                    �?      �?             @@�       �                    �M@�IєX�?
             1@�       �                    �?r�q��?             @������������������������       �                      @�       �       	             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �        	             .@�       �                    @E@�G\�c�?)            @P@������������������������       �                     $@�       �                    �?D7�J��?#            �K@�       �       	          ����?\�Uo��?             C@�       �                    @L@�!���?             A@�       �                    �?������?             >@������������������������       �                     .@�       �       
             �?��S���?             .@������������������������       �                      @�       �                   Pd@��
ц��?             *@�       �                    �?���|���?	             &@�       �                    �?�z�G��?             $@�       �                   @q@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   c@      �?             @������������������������       �                      @�       �                   p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @�t����?             1@�       �       	          @33�?z�G�z�?             .@������������������������       �                     &@�       �                    �N@      �?             @�       �                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?�8=�?           �y@�       �                    �?68��1��?N            �^@�       �                   �`@F�����?8            �V@�       �                   �U@ףp=
�?             >@������������������������       �                     �?�       �                   `]@ 	��p�?             =@������������������������       �                     0@�       �                   �^@8�Z$���?             *@������������������������       �                      @������������������������       �                     &@�       �                   `T@�������?'             N@������������������������       �                     *@�       �       	          ����?֭��F?�?             �G@�       �                    �?�!���?             A@�       �                   �d@؇���X�?             @������������������������       �                     @�       �                    �H@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��}*_��?             ;@�       �                   �b@�n_Y�K�?             :@�       �                     N@���N8�?             5@�       �                    ]@z�G�z�?             4@�       �                   d@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �K@��S�ۿ?             .@������������������������       �                     (@�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �?��
ц��?	             *@�       �       	          ����?���|���?             &@������������������������       �                     @�       �                   @_@�q�q�?             @�       �                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                   Pd@     ��?             @@�       �       	          ����?д>��C�?             =@�       �                    �?�n_Y�K�?             *@�       �                   P`@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   �Z@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     0@�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   @c@DK{22�?�             r@�       �                    �N@�û��|�?             7@�       �                   �b@��S���?
             .@�       �       	          `ff�?��
ц��?	             *@������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �_@      �?              @�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�             	             @ p�/��?�            �p@�                         �g@�zvܰ?�            �p@�       �                    @L@������?�            Pp@�       �                   @[@@f��F�?~             i@�       �                   �Z@�8��8��?	             (@������������������������       �                     $@�       �                   �o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        u            �g@�       �                    �?ףp=
�?"             N@������������������������       �                     >@�                          @z�G�z�?             >@�                          �?�8��8��?             8@�       �                   pa@�KM�]�?             3@������������������������       �                     @�       �                    �L@r�q��?             (@������������������������       �                     �?�                          ps@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     @                          O@�q�q�?             @������������������������       �                     @������������������������       �                      @                         d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM	KK��h_�B�       @z@      @      V@      z@     �F@     �u@      7@     �q@      �?     �T@      �?      3@              3@      �?                     �O@      6@      i@      &@     �K@      @       @               @      @              @     �J@      @     �J@              .@      @      C@              5@      @      1@              @      @      *@      @      @      @      @      �?               @      @       @      @      �?      @              @      �?      �?              �?      �?              �?                       @       @                      @       @              &@      b@              B@      &@     @[@      $@     @P@      @      @              @      @              @      N@      @      L@      �?      @      �?                      @       @      J@      �?     �I@      �?      @              @      �?       @      �?                       @              G@      �?      �?      �?                      �?      @      @      �?              @      @      @                      @      �?      F@      �?      *@              @      �?      "@      �?      �?      �?                      �?               @              ?@      6@     �P@      $@      K@      @     �J@      @     �J@      @      B@      @      A@      @      .@      �?      *@      �?       @      �?       @              �?      �?      �?              �?      �?                      @              @       @       @       @                       @              3@       @       @       @                       @              1@       @              @      �?              �?      @              (@      (@      &@      @      @              @      @      @      @      @      @              @      @      �?      @                      �?       @                      �?      �?      @              @      �?      �?      �?                      �?     �E@     �Q@      @     �E@      @      (@      @      �?      @                      �?              &@      �?      ?@      �?      0@      �?      @               @      �?      @              @      �?                      &@              .@      C@      ;@      $@              <@      ;@      7@      .@      7@      &@      6@       @      .@              @       @               @      @      @      @      @      @      @      @      �?      @                      �?               @              �?               @      �?      @               @      �?      �?      �?                      �?              @      @      (@      @      (@              &@      @      �?      �?      �?              �?      �?               @               @             �t@      T@     �O@     �M@      L@      A@      ;@      @              �?      ;@       @      0@              &@       @               @      &@              =@      ?@              *@      =@      2@      7@      &@      @      �?      @              �?      �?      �?                      �?      1@      $@      0@      $@      0@      @      0@      @       @      @              @       @              ,@      �?      (@               @      �?       @                      �?              �?              @      �?              @      @      @      @              @      @       @      �?       @      �?                       @      @               @              @      9@      @      8@      @       @      �?      @      �?                      @      @       @               @      @                      0@       @      �?       @                      �?     �p@      5@      ,@      "@      @       @      @      @      @                      @               @      @      �?       @      �?       @                      �?      @             �o@      (@     �o@      "@     �o@      @      i@      �?      &@      �?      $@              �?      �?              �?      �?             �g@              K@      @      >@              8@      @      6@       @      1@       @      @              $@       @              �?      $@      �?      $@                      �?      @               @      @              @       @              �?       @      �?                       @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���yhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM!hwh(h+K ��h-��R�(KM!��h~�B8?         |                    @K@�$�����?P           ��@       C                    �?�"����?0           ~@              
             �?�|ew���?�             k@                          �i@��*��?]            `a@                           �D@(;L]n�?(             N@                           b@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?	       
                   �U@@��8��?              H@������������������������       �                     �?������������������������       �                    �G@              	          ����?���!���?5            �S@                           �?4�2%ޑ�?            �A@                           �C@      �?             $@������������������������       �                      @              	          ����?      �?              @������������������������       �                      @                          �b@r�q��?             @������������������������       �                     @������������������������       �                     �?                           `@H%u��?             9@������������������������       �                     ,@                           �F@���!pc�?             &@������������������������       �                      @������������������������       �                     @                          �a@`���i��?             F@������������������������       �                     E@                          �m@      �?              @������������������������       �                     �?������������������������       �                     �?       2                   �_@��c�%�?.            @S@        %                   �g@�xGZ���?            �A@!       "                    �?      �?             0@������������������������       �                     (@#       $                   �X@      �?             @������������������������       �                      @������������������������       �                      @&       1                   �^@�d�����?             3@'       *                    @F@@�0�!��?             1@(       )                   �q@      �?             @������������������������       �                      @������������������������       �                      @+       0                    �?$�q-�?             *@,       /                    �G@      �?              @-       .                    �F@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @3       8                   �b@��s����?             E@4       5       	          433�? ��WV�?             :@������������������������       �                     7@6       7                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @9       >                    �?     ��?             0@:       =                   �b@�z�G��?             $@;       <       	          `ffֿ      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @?       B       	             �?�q�q�?             @@       A                   (p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @D       O                   �c@��c��?�            �p@E       J                     G@���N8�?             5@F       I                    @      �?              @G       H                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @K       N       
             �?$�q-�?             *@L       M                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@P       ]                    �?����B��?�            �n@Q       R                    @H@���N8�?5             U@������������������������       �                    �E@S       T                   �Z@������?            �D@������������������������       �                      @U       V                    g@�7��?            �C@������������������������       �                     �?W       X                   @a@P�Lt�<�?             C@������������������������       �                     :@Y       Z                    �?�8��8��?             (@������������������������       �                     $@[       \                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?^       i       	          ����?ףp=��?b             d@_       h       
             �?PF��t<�?L            �_@`       a                   ``@�q�q�?	             (@������������������������       �                     �?b       e       	          ����?���!pc�?             &@c       d                     C@      �?              @������������������������       �                     �?������������������������       �                     @f       g       	          pff�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        C            �\@j       k                    �?�eP*L��?            �@@������������������������       �                     @l       {                    �?X�<ݚ�?             ;@m       z       
             �?�LQ�1	�?             7@n       w       	          ����?�X����?             6@o       v                   �e@��
ц��?	             *@p       u                   �l@�q�q�?             (@q       t                   �h@r�q��?             @r       s                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?x       y       
             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @}       �                    �?,y)�S�?            P{@~       �                    �?P�TΧ��?�            �p@       �                    �?h�x�P��?o             e@�       �                   �a@�eP*L��?$            �K@�       �                   @Z@z�J��?            �G@������������������������       �                      @�       �                   �c@�ݏ^���?            �F@�       �                   @E@D^��#��?            �D@�       �                   `]@�C��2(�?             &@������������������������       �                     @�       �       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                     P@�z�G��?             >@�       �                    @N@؇���X�?             5@�       �       
             �?�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     &@�       �                    �?�q�q�?             "@������������������������       �                      @�       �                   0b@؇���X�?             @������������������������       �                     @�       �       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   0l@      �?              @������������������������       �                     @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @N@����?K            @\@�       �                    �?�z�6�?'             O@������������������������       �                     2@�       �                   Pd@v�X��?             F@�       �       	          ����?^����?            �E@�       �       
             �?�q�q�?             (@������������������������       �                     �?�       �                     L@���!pc�?             &@������������������������       �                      @�       �                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �       
             �?��� ��?             ?@������������������������       �                     :@�       �                   �\@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    �?�IєX�?$            �I@�       �                   �q@z�G�z�?             $@������������������������       �                     @�       �                   0a@�q�q�?             @������������������������       �                     �?�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   ``@��Y��]�?            �D@�       �                   p@      �?
             0@������������������������       �                     (@�       �                   �p@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     9@�       �                   �[@@9G��??            �X@������������������������       �                     D@�       �                    �? 	��p�?(             M@������������������������       �                     @�       �                   x@�:�]��?#            �I@�       �                    �R@@9G��?"            �H@������������������������       �        !            �G@������������������������       �                      @������������������������       �                      @�       �                   �d@�\��N��?r            `e@�       �       
             �?�������?             A@�       �                   �c@�LQ�1	�?             7@�       �                    �?�����?             5@�       �       	          hff@      �?              @�       �                    �?�q�q�?             @�       �                   �]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �        	             *@�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     Q@�eP*L��?             &@�       �                    �?؇���X�?             @������������������������       �                     @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�             
             �?���5��?Z             a@�       �                    �?�q�q�?1             R@�       �                    �?z�G�z�?             $@�       �                    �?�����H�?             "@�       �                    @L@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �[@r֛w���?)             O@������������������������       �                     @�       �       
             �?V�a�� �?'             M@�       �                   �^@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �a@���c���?$             J@�       �                    @      �?             @@�       �                   �`@(;L]n�?             >@�       �                   �r@؇���X�?             @������������������������       �                     @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@�       �                   c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   b@      �?             4@������������������������       �                      @�                          �?r�q��?             2@�       �                    �L@      �?
             (@������������������������       �                     �?�       �       	          pff�?"pc�
�?	             &@������������������������       �                     �?�                          �O@ףp=
�?             $@             	          033@z�G�z�?             @                        @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @             	             @�?�<��?)            @P@                         �?     ��?(             P@	                         @M@V�a�� �?             =@
                         �?�q�q�?             2@            	          @33�?���Q��?             @                        Hv@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                        @_@�	j*D�?	             *@            	          pff�?      �?             @������������������������       �                     @������������������������       �                     �?                         @L@�����H�?             "@������������������������       �                     @                         c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@                        �c@��?^�k�?            �A@������������������������       �                     :@                         �N@�����H�?             "@������������������������       �                     @                        �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�t�b�     h�h(h+K ��h-��R�(KM!KK��h_�B       `z@      @     �q@     @h@     �N@     `c@      &@      `@       @      M@      �?      &@              &@      �?              �?     �G@      �?                     �G@      "@     �Q@       @      ;@      @      @               @      @      @               @      @      �?      @                      �?      @      6@              ,@      @       @               @      @              �?     �E@              E@      �?      �?      �?                      �?      I@      ;@      0@      3@       @      ,@              (@       @       @               @       @              ,@      @      ,@      @       @       @       @                       @      (@      �?      @      �?      @      �?      @                      �?      @              @                       @      A@       @      9@      �?      7@               @      �?              �?       @              "@      @      @      @      @      �?              �?      @                       @       @      @       @      �?              �?       @                      @     @l@     �C@      @      0@      @      @      @       @               @      @                       @      �?      (@      �?       @      �?                       @              $@     �k@      7@      T@      @     �E@             �B@      @               @     �B@       @              �?     �B@      �?      :@              &@      �?      $@              �?      �?              �?      �?             �a@      3@     �^@      @       @      @              �?       @      @      @      �?              �?      @              �?       @               @      �?             �\@              2@      .@      @              (@      .@       @      .@      @      .@      @      @      @      @      @      �?      �?      �?      �?                      �?      @                      @      �?              �?       @      �?                       @      �?              @             �`@     �r@     �F@     �k@     �D@     �_@      9@      >@      8@      7@       @              6@      7@      6@      3@      �?      $@              @      �?      @      �?                      @      5@      "@      2@      @      @      @              @      @              &@              @      @       @              �?      @              @      �?       @      �?                       @              @      �?      @              @      �?      �?      �?                      �?      0@     @X@      *@     �H@              2@      *@      ?@      (@      ?@       @      @              �?       @      @       @              @      @              @      @              @      ;@              :@      @      �?      @                      �?      �?              @      H@       @       @              @       @      �?      �?              �?      �?              �?      �?              �?      D@      �?      .@              (@      �?      @      �?                      @              9@      @     �W@              D@      @      K@              @      @     �G@       @     �G@             �G@       @               @             �V@     @T@      "@      9@      @      4@       @      3@       @      @       @      @       @       @       @                       @               @               @              *@      �?      �?      �?                      �?      @      @      @      �?      @              �?      �?              �?      �?                      @     @T@      L@      8@      H@       @       @       @      �?      @      �?      @                      �?      @                      �?      0@      G@      @              (@      G@      @      �?              �?      @              @     �F@       @      >@      �?      =@      �?      @              @      �?      �?              �?      �?                      7@      �?      �?              �?      �?              @      .@       @              @      .@      @      "@      �?               @      "@      �?              �?      "@      �?      @      �?      �?              �?      �?                      @              @              @     �L@       @     �L@      @      7@      @      (@      @      @       @      �?       @               @      �?               @              "@      @      �?      @              @      �?               @      �?      @               @      �?       @                      �?      &@              A@      �?      :@               @      �?      @              �?      �?              �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���3hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK݅�h~�BX0         �       
             �?2���xA�?;           ��@       %                    �?��USa�?G           ��@       "                   �c@���Q��?0             T@       !                    �?�&�5y�?&             O@                           �O@�&!��?            �E@              	          ����?<ݚ)�?             B@                          �_@�q�q�?             8@                          Pf@�����H�?             "@	       
                    �D@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           @H@���Q��?
             .@������������������������       �                     @                          `^@      �?              @                           �?�q�q�?             @������������������������       �                     �?                          xu@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          �`@�8��8��?	             (@                           �I@      �?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �?؇���X�?             @������������������������       �                     @               	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             3@#       $                    �?r�q��?
             2@������������������������       �                     @������������������������       �                     .@&       Y                    �?l�$֧X�?           0|@'       .                   i@ �tI���?�            �t@(       )                   �_@�[�mT�?V            �a@������������������������       �        7            �V@*       +                   pb@p���?             I@������������������������       �                     C@,       -                    �G@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@/       L                    �?��Y���?w            �g@0       K                    @M@�2c�$��?Z             b@1       2                   �S@�8�l��?B            �Z@������������������������       �                     �?3       4                   �Z@ >�֕�?A            @Z@������������������������       �                     �?5       J       	          ����?��s�n�?@             Z@6       G                    @L@85�}C�?&            �N@7       8                    �?h�����?#             L@������������������������       �                     "@9       F                   �`@`�q�0ܴ?            �G@:       C                   ``@ 	��p�?             =@;       <                    �? 7���B�?             ;@������������������������       �                     @=       B                    \@���N8�?             5@>       ?                   �Z@�����H�?             "@������������������������       �                     @@       A                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             (@D       E                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             2@H       I                   ``@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                    �E@������������������������       �                    �C@M       X       	             �?�㙢�c�?             G@N       Q                    Y@��.k���?	             1@O       P                   (q@؇���X�?             @������������������������       �                     @������������������������       �                     �?R       S       	             �?z�G�z�?             $@������������������������       �                     @T       U                    `@      �?             @������������������������       �                     �?V       W                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     =@Z       w                   P`@������?J             ^@[       t                   0f@�d�K���?)            �P@\       _                    @E@T����1�?$             M@]       ^                   o@r�q��?             @������������������������       �                     @������������������������       �                     �?`       o                   �n@R�}e�.�?             J@a       n                   �m@�q�q�?             B@b       e                    Y@���!pc�?            �@@c       d                    X@      �?              @������������������������       �                     @������������������������       �                     @f       g                    `@�J�4�?             9@������������������������       �                     3@h       m                    @�q�q�?             @i       j                   @`@z�G�z�?             @������������������������       �                      @k       l                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @p       s                    �?      �?	             0@q       r                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     (@u       v       	          033@�����H�?             "@������������������������       �                      @������������������������       �                     �?x       �                    @0��_��?!            �J@y       z                   `b@`Ӹ����?            �F@������������������������       �                     9@{       �                    �Q@ףp=
�?             4@|       }                    @N@�}�+r��?
             3@������������������������       �                     .@~                           �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   l@      �?              @������������������������       �                     @�       �       
             �?���Q��?             @������������������������       �                      @�       �                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    I@J3�xH��?�            0x@�       �       	            �?��2(&�?             F@�       �                   a@������?
             1@�       �       	          033�؇���X�?             ,@������������������������       �                     @�       �       	             п�<ݚ�?             "@������������������������       �                     �?�       �       	          ����?      �?              @�       �                   �\@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   0d@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    c@�>����?             ;@�       �                    �M@ �q�q�?             8@������������������������       �                     0@�       �       	          `ff�?      �?              @������������������������       �                     @�       �                    a@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�x=Fh_�?�            pu@�       �                    �?b�2�tk�?9            �V@�       �                   �q@����X�?            �A@�       �       	          ����?�G��l��?             5@�       �                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                    m@"pc�
�?             &@�       �                   �j@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     ,@�       �                    �?"pc�
�?&            �K@�       �       	          033�?�C��2(�?             F@�       �                   pf@Du9iH��?            �E@�       �                    Z@�(\����?             D@������������������������       �                     �?������������������������       �                    �C@�       �                    �B@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    @M@�eP*L��?
             &@�       �                    �?�q�q�?             @�       �       	          ����?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �       	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �`@0��kS֣?�            �o@�       �                    @L@�������?h            �d@������������������������       �        `             c@�       �                   �p@$�q-�?             *@�       �                   �a@r�q��?             @������������������������       �                     @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @`��F:u�?5            �U@�       �                    a@F|/ߨ�?1            @T@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �c@�(�Tw�?/            �S@�       �       	          ����?P�Lt�<�?             C@�       �                    �?`2U0*��?             9@������������������������       �                      @�       �                   @c@�nkK�?             7@������������������������       �                     6@������������������������       �                     �?������������������������       �        	             *@������������������������       �                     D@�       �                   �a@�q�q�?             @������������������������       �                     @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       Px@     ��@      T@     0|@      @@      H@      1@     �F@      1@      :@      &@      9@      $@      ,@      �?       @      �?       @               @      �?                      @      "@      @      @               @      @       @      �?      �?              �?      �?      �?                      �?              @      �?      &@      �?      @      �?      �?              �?      �?                       @               @      @      �?      @              @      �?              �?      @                      3@      .@      @              @      .@              H@     0y@      0@     �s@      �?     `a@             �V@      �?     �H@              C@      �?      &@      �?                      &@      .@      f@      @     @a@      @     �X@      �?              @     �X@      �?              @     �X@      @      L@       @      K@              "@       @     �F@       @      ;@      �?      :@              @      �?      4@      �?       @              @      �?       @               @      �?                      (@      �?      �?      �?                      �?              2@      @       @      @                       @             �E@             �C@       @      C@       @      "@      @      �?      @                      �?       @       @              @       @       @      �?              �?       @               @      �?                      =@      @@      V@      ;@      D@      3@     �C@      @      �?      @                      �?      ,@      C@      (@      8@      "@      8@      @      @              @      @              @      5@              3@      @       @      @      �?       @               @      �?              �?       @                      �?      @               @      ,@       @       @       @                       @              (@       @      �?       @                      �?      @      H@       @     �E@              9@       @      2@      �?      2@              .@      �?      @              @      �?              �?              @      @              @      @       @       @              �?       @               @      �?             Ps@     �S@      @      C@      @      *@       @      (@              @       @      @      �?              �?      @      �?      @      �?                      @              �?       @      �?       @                      �?       @      9@      �?      7@              0@      �?      @              @      �?      @      �?                      @      �?       @      �?                       @     �r@      D@     �K@     �A@      $@      9@      $@      &@       @       @       @                       @       @      "@       @      @              @       @                      @              ,@     �F@      $@      D@      @      D@      @     �C@      �?              �?     �C@              �?       @      �?                       @              �?      @      @      @       @      @       @      @                       @      �?              �?      @      �?                      @      o@      @     �d@      �?      c@              (@      �?      @      �?      @              �?      �?              �?      �?              @             �T@      @     �S@       @       @      �?              �?       @             @S@      �?     �B@      �?      8@      �?       @              6@      �?      6@                      �?      *@              D@              @       @      @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��4hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�5         �       
             �?�LT ���?E           ��@       K                    �?
�GN��?N           ��@                           �?l��\��?�            `w@              	          ����?��]�T��?            �D@                          c@     ��?             0@                          �j@8�Z$���?	             *@                            H@�q�q�?             @������������������������       �                     �?	       
                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     @                          h@�J�4�?             9@                           �?���Q��?             @������������������������       �                      @������������������������       �                     @                          �_@ףp=
�?             4@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �        
             ,@                          `R@@-�_ .�?�            �t@                           a@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           Z@�6,r➷?�            �t@                          �Y@z�G�z�?             .@������������������������       �                     (@������������������������       �                     @       J                   �e@H�C.B�?�            �s@        !       	          ����?��j��Ѳ?�            �s@������������������������       �        )            @Q@"       '       	          ����?(z�Iiٷ?�            �n@#       $                    @M@և���X�?             @������������������������       �                     @%       &                   �_@      �?             @������������������������       �                     �?������������������������       �                     @(       ?                    �?0x�!���?�            �m@)       <                    �R@ _�@�Y�?l            �e@*       ;                    �?��f�{��?j            �e@+       ,                    �? ������?L            �_@������������������������       �                    �@@-       .                   �d@����D��?7            @W@������������������������       �                     ;@/       0                   @a@Pa�	�?*            �P@������������������������       �                    �@@1       2                    �?�FVQ&�?            �@@������������������������       �                     @3       4                   �f@@4և���?             <@������������������������       �                     �?5       6       
             �? 7���B�?             ;@������������������������       �                     @7       8                   �p@�nkK�?             7@������������������������       �                     3@9       :                   �q@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     G@=       >                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?@       E                   �_@     p�?(             P@A       B                    @J@և���X�?             @������������������������       �                     �?C       D                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     @F       I       	             �?0�)AU��?#            �L@G       H                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        !             K@������������������������       �                     �?L       �                    �?i����?d            @c@M       b                   a@�p ��?P            �^@N       [                   pm@��Hg���?            �F@O       V                     P@J�8���?             =@P       U                    �?@4և���?	             ,@Q       T                   �Z@      �?              @R       S                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @W       X                    �?���Q��?	             .@������������������������       �                      @Y       Z                   �k@؇���X�?             @������������������������       �                     @������������������������       �                     �?\       ]       	             �?      �?             0@������������������������       �                     "@^       _                   �r@؇���X�?             @������������������������       �                     @`       a                    �?      �?              @������������������������       �                     �?������������������������       �                     �?c       �                   �e@�q�q�?3            �S@d       e       
             �?      �?+             P@������������������������       �                     @f                           �?6�iL�?(            �M@g       h                    �F@�GN�z�?             F@������������������������       �                     ,@i       j                   �g@�q�q�?             >@������������������������       �                     @k       l                     H@������?             ;@������������������������       �                      @m       r                   �b@z�G�z�?             9@n       o       	          833�?���Q��?             @������������������������       �                      @p       q                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @s       x                    �L@R���Q�?             4@t       w       	          `ff�?$�q-�?
             *@u       v                   @a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@y       z                    �?����X�?             @������������������������       �                     �?{       ~                   �x@r�q��?             @|       }                    �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   (p@���Q��?
             .@�       �                   b@ףp=
�?             $@������������������������       �                     @�       �                   @`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   g@����X�?             ,@�       �                   f@r�q��?             (@������������������������       �                     @�       �                   �p@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                   `c@�n`���?             ?@�       �       	          ����?\-��p�?             =@�       �                    �?�<ݚ�?             2@�       �                    �?�	j*D�?	             *@�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �Z@z�G�z�?             $@�       �                   `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     &@������������������������       �                      @�       �                    �?f�ȭ��?�            `x@�       �                    �?����3�?�             t@�       �       	            �?�	j*D�?L            @]@�       �                   pc@��f��?6            @V@�       �                   @_@��<b�ƥ?             G@�       �                    @P@      �?             0@������������������������       �                     .@������������������������       �                     �?������������������������       �                     >@�       �                   �f@�&!��?            �E@�       �                    b@��
P��?            �A@�       �                    �?�P�*�?             ?@������������������������       �                     "@�       �                    �?8�A�0��?             6@������������������������       �                     @�       �                    @G@���Q��?	             .@������������������������       �                      @�       �                   �d@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �u@X�Cc�?             <@�       �                    �C@      �?             8@������������������������       �                     �?�       �                   0c@��<b���?             7@�       �       	             �?؇���X�?             5@�       �                    �M@@4և���?
             ,@������������������������       �                     "@�       �                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?����X�?             @�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?z�G�z�?             @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    @L@�<e3�?�            �i@�       �                   �g@�C��2(�?p             f@�       �                    �?���ib#�?o            �e@�       �                   @`@���7�?             6@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     3@�       �                    �?��ꤘ�?`             c@������������������������       �        O             `@�       �                    T@`2U0*��?             9@�       �                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     6@������������������������       �                     �?�       �                    �?д>��C�?             =@������������������������       �                     $@�       �                   ps@�d�����?             3@�       �                    �M@@�0�!��?             1@�       �                    d@      �?              @������������������������       �                     @�       �                   �a@      �?             @������������������������       �                      @�       �                    i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                      @�       �                   pc@�������?&             Q@�       �                   �Y@�I�w�"�?             C@������������������������       �                      @�       �                    �?tk~X��?             B@�       �                   Xv@HP�s��?             9@�       �                    �? �q�q�?             8@������������������������       �        
             3@�       �                   `\@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                    V@�eP*L��?             &@������������������������       �                     @������������������������       �                     @�       �                    �?z�G�z�?             >@������������������������       �                     @������������������������       �                     8@�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       �y@     �@     �Y@     �z@     �@@     Pu@      .@      :@      &@      @      &@       @      �?       @              �?      �?      �?      �?                      �?      $@                      @      @      5@       @      @       @                      @       @      2@       @      @       @                      @              ,@      2@     �s@       @      �?       @                      �?      0@     �s@      @      (@              (@      @              *@     �r@      (@     �r@             @Q@      (@      m@      @      @      @              �?      @      �?                      @       @     �l@      @     `e@       @     @e@       @      _@             �@@       @     �V@              ;@       @      P@             �@@       @      ?@              @       @      :@      �?              �?      :@              @      �?      6@              3@      �?      @      �?                      @              G@      �?      �?              �?      �?              @     �M@      @      @              �?      @       @               @      @              �?      L@      �?       @      �?                       @              K@      �?             @Q@     @U@     �O@      N@      &@      A@      $@      3@      �?      *@      �?      @      �?      �?      �?                      �?              @              @      "@      @       @              �?      @              @      �?              �?      .@              "@      �?      @              @      �?      �?      �?                      �?      J@      :@      H@      0@      @             �E@      0@      A@      $@      ,@              4@      $@              @      4@      @               @      4@      @      @       @       @              �?       @      �?                       @      1@      @      (@      �?       @      �?       @                      �?      $@              @       @              �?      @      �?       @      �?              �?       @              @              "@      @      "@      �?      @              @      �?      @                      �?              @      @      $@       @      $@              @       @      @              @       @               @              @      9@      @      9@      @      ,@      @      "@       @      �?              �?       @               @       @       @      �?              �?       @                      @              @              &@       @             ps@     �S@     `q@      F@     @T@      B@     �Q@      2@     �F@      �?      .@      �?      .@                      �?      >@              :@      1@      2@      1@      2@      *@      "@              "@      *@              @      "@      @       @              �?      @              @      �?                      @       @              $@      2@      @      2@      �?              @      2@      @      2@      �?      *@              "@      �?      @              @      �?               @      @      �?      �?              �?      �?              �?      @      �?      �?      �?                      �?              @       @              @             �h@       @     �e@      @     �e@       @      5@      �?       @      �?       @                      �?      3@              c@      �?      `@              8@      �?       @      �?       @                      �?      6@                      �?      8@      @      $@              ,@      @      ,@      @      @      @      @              �?      @               @      �?      �?      �?                      �?      "@                       @     �@@     �A@      "@      =@       @              @      =@       @      7@      �?      7@              3@      �?      @              @      �?              �?              @      @              @      @              8@      @              @      8@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���
hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK녔h~�Bh3         �                    �?x��X���?Z           ��@       M       
             �?&\@��??           p@       B                   �a@�h����?�            pw@              	          833�?���x��?�            �n@������������������������       �        $            �J@                          0h@�q�Q�?y             h@                           �?�8���?"             M@                           �Q@��a�n`�?             ?@	       
                    �?XB���?             =@������������������������       �        
             3@              
             �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                      @������������������������       �                     ;@       ?                    �?V�L��?W            �`@                           �?��U/��?H            �\@              	          ����?���!pc�?             6@                          �a@�r����?
             .@              	          ����?�<ݚ�?             "@������������������������       �                     �?                          a@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                           �?և���X�?             @                           �O@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       *                    @J@�3Ea�$�?9             W@        %                    �?ףp=
�?             >@!       $                    �F@����X�?             @"       #                    ]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @&       )                   �j@�nkK�?             7@'       (                     D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     5@+       ,                    �J@j�g�y�?%             O@������������������������       �                     @-       >                   �b@&y�X���?$             M@.       7                    �L@H�ՠ&��?!             K@/       6       	             �?����X�?             5@0       1                    ^@�q�q�?             "@������������������������       �                      @2       3                   `W@և���X�?             @������������������������       �                      @4       5                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@8       9                    `@Pa�	�?            �@@������������������������       �                     3@:       =                    �?@4և���?
             ,@;       <                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                     @@       A                   �S@P���Q�?             4@������������������������       �                     �?������������������������       �                     3@C       L       	          ����?0�ޤ��?N            @`@D       K                    �H@Hn�.P��?'             O@E       J                    �?և���X�?             @F       G                    �D@���Q��?             @������������������������       �                      @H       I                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        "            �K@������������������������       �        '             Q@N       w                    �?     ��?T             `@O       h       	          ����?6n�
$)�?>            �W@P       W                   �b@��<b���?,            @Q@Q       V                    �?�?�|�?            �B@R       S       	            �?XB���?             =@������������������������       �                     :@T       U                    V@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @X       ]                   �_@     ��?             @@Y       Z                   `i@z�G�z�?             $@������������������������       �                     @[       \                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     @^       c                    �?���!pc�?             6@_       b                     N@@�0�!��?	             1@`       a                   @b@      �?             0@������������������������       �                     ,@������������������������       �                      @������������������������       �                     �?d       e                   @`@���Q��?             @������������������������       �                      @f       g                    h@�q�q�?             @������������������������       �                     �?������������������������       �                      @i       l                    �F@ �o_��?             9@j       k                   0b@      �?             @������������������������       �                     �?������������������������       �                     @m       v                    c@��s����?             5@n       u                    @N@�KM�]�?             3@o       p       	          pff�?�<ݚ�?             "@������������������������       �                     �?q       r       	             �?      �?              @������������������������       �                     @s       t                   ``@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                      @x       }                   ``@@�0�!��?             A@y       |                    �?���N8�?             5@z       {                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     2@~                           �I@�n_Y�K�?             *@������������������������       �                     @�       �       	          ����?�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       
             �?Ԡ��	�?           �y@�       �                   �o@�F}ʽx�?n            �b@�       �                   �`@༉p���?M            �Z@�       �                    �?�p ��?            �D@������������������������       �                     �?�       �                    �?      �?             D@�       �                   @j@���Q��?             @�       �       	          `ff�?      �?             @�       �                   `Y@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   �^@ >�֕�?            �A@�       �       	             �?8�Z$���?
             *@�       �       	          ���ٿ�<ݚ�?             "@������������������������       �                     �?�       �                   `]@      �?              @������������������������       �                     @�       �                    V@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     6@�       �                   0g@:ɨ��?/            �P@�       �                    �G@և���X�?
             ,@������������������������       �                     @�       �                    �?���!pc�?             &@������������������������       �                     @�       �       	             @      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @L@�θ�?%             J@�       �                    �?�S����?             C@������������������������       �        
             *@�       �                    �F@�+e�X�?             9@�       �                   �l@$�q-�?             *@������������������������       �                     $@�       �                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �m@�q�q�?             (@�       �                   �d@�z�G��?             $@�       �                    �H@      �?              @�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �       	          ����?և���X�?             ,@������������������������       �                     @�       �                    @���!pc�?	             &@�       �                   �b@և���X�?             @������������������������       �                     @�       �                    [@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?fP*L��?!             F@�       �                     L@���Q��?
             $@������������������������       �                      @�       �                   �a@      �?              @������������������������       �                     @�       �                   pb@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?l��\��?             A@�       �                    �?@�0�!��?             1@�       �                   �b@d}h���?             ,@�       �                   �r@8�Z$���?
             *@������������������������       �                     $@�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        	             1@�       �                   �O@���7�?�            �p@�       �       	          ����?      �?             $@������������������������       �                     @������������������������       �                     @�       �                   �g@���Wq�?�            �o@�       �       	             @@7���?�            `o@�       �                   �b@@Lb�G�?�            @o@������������������������       �        G            �\@�       �                   �s@����?�?\            �`@�       �                   �d@ ���z��?U            �_@�       �                    �?`'�J�?!            �I@�       �                    @L@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     G@������������������������       �        4             S@�       �                    �?      �?              @�       �                    w@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       0z@     0@      [@     �x@     �D@     �t@      C@     �i@             �J@      C@     @c@      @     �K@      @      <@      �?      <@              3@      �?      "@      �?                      "@       @                      ;@     �A@     �X@      A@      T@      0@      @      *@       @      @       @              �?      @      �?      @                      �?      @              @      @      @      �?              �?      @                      @      2@     �R@      @      ;@       @      @       @       @       @                       @              @      �?      6@      �?      �?              �?      �?                      5@      .@     �G@      @              &@     �G@      @     �G@      @      .@      @      @       @              @      @               @      @      �?              �?      @                      (@      �?      @@              3@      �?      *@      �?       @               @      �?                      &@      @              �?      3@      �?                      3@      @     �_@      @     �M@      @      @      @       @       @              �?       @      �?                       @               @             �K@              Q@     �P@     �N@     �N@     �@@      K@      .@      B@      �?      <@      �?      :@               @      �?              �?       @               @              2@      ,@       @       @              @       @      @       @                      @      0@      @      ,@      @      ,@       @      ,@                       @              �?       @      @               @       @      �?              �?       @              @      2@      @      �?              �?      @              @      1@       @      1@       @      @      �?              �?      @              @      �?      �?      �?                      �?              $@       @              @      <@      �?      4@      �?       @      �?                       @              2@      @       @      @              �?       @      �?                       @     ps@      Z@     �M@      W@      J@     �K@      @     �A@      �?              @     �A@      @       @      @      �?       @      �?              �?       @              �?                      �?       @     �@@       @      &@       @      @              �?       @      @              @       @       @               @       @                      @              6@      G@      4@      @       @      @              @       @              @      @      �?       @              �?      �?              �?      �?              D@      (@      @@      @      *@              3@      @      (@      �?      $@               @      �?              �?       @              @      @      @      @      @      �?       @      �?              �?       @              @                       @               @       @      @              @       @      @      @      @      @              �?      @      �?                      @      @              @     �B@      @      @       @               @      @              @       @       @      �?              �?       @      �?                       @      @      ?@      @      ,@      @      &@       @      &@              $@       @      �?              �?       @              �?                      @              1@     �o@      (@      @      @      @                      @     �n@      @     �n@      @     �n@      @     �\@             �`@      @     @_@       @     �H@       @      @       @      @                       @      G@              S@              @      �?      �?      �?              �?      �?              @                      �?              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJI�whG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �                    �?X�<ݚ�?N           ��@       M       
             �?��<b���?<           0~@       *       	             �?�d�S��?�            �u@       %                    �?�S�w���?m            `d@                          @l@�s�n_�?G             Z@                           �?��<b�ƥ?!             G@������������������������       �                     ?@                          �X@��S�ۿ?	             .@	       
       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@       "                   `a@�f7�z�?&             M@              	          ����?�s��:��?             C@                          �b@�����H�?             "@������������������������       �                     @                          �p@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?8^s]e�?             =@                           @I@�C��2(�?             &@                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                           `@X�<ݚ�?             2@                           `P@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @       !                   �r@�q�q�?             "@                           `Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @#       $                   �l@R���Q�?             4@������������������������       �                     @������������������������       �        
             1@&       '                   Pz@���#�İ?&            �M@������������������������       �        $             L@(       )       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?+       ,                   �U@P��a4�?v            �g@������������������������       �                     @-       4                   @^@x�û��?u             g@.       3                    �J@�E�����?6            �V@/       2                   �_@P���Q�?             4@0       1       	             @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             ,@������������������������       �        (            �Q@5       :                   @\@=QcG��??            �W@6       9                   �k@�z�G��?             $@7       8                   �X@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @;       >                   �^@h�����?7             U@<       =                     N@؇���X�?             @������������������������       �                     @������������������������       �                     �??       F                   �g@�g<a�?2            @S@@       E                    @J@$�q-�?	             *@A       B                    �?      �?             @������������������������       �                      @C       D       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@G       H                    @M@     ��?)             P@������������������������       �                     A@I       L                   �a@(;L]n�?             >@J       K                    �M@@4և���?	             ,@������������������������       �                     �?������������������������       �                     *@������������������������       �                     0@N       w       	          ����?��e���?Y            �`@O       T                   �X@��Sݭg�?9            �S@P       S                   �V@����X�?             @Q       R       	             ��q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @U       j                    �M@@���?T�?4            �Q@V       a                   �_@t�6Z���?(            �K@W       X                   �b@�����?             3@������������������������       �                     $@Y       `                    �I@�q�q�?             "@Z       _                    �?���Q��?             @[       \                    �?      �?             @������������������������       �                     �?]       ^                    \@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @b       c       	          `ffֿ�X�<ݺ?             B@������������������������       �                     �?d       e                    �?��?^�k�?            �A@������������������������       �                     @f       i                    �D@h�����?             <@g       h                   @b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     9@k       v       	          ����?     ��?             0@l       o                    _@���|���?	             &@m       n                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?p       q                    �?      �?              @������������������������       �                     @r       u                   @b@�q�q�?             @s       t                     P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @x       �                   0e@r�q��?              K@y       ~                    �?�t����?            �I@z       {                    [@z�G�z�?             4@������������������������       �                     �?|       }                   �`@�S����?             3@������������������������       �        	             0@������������������������       �                     @       �                    �?`Jj��?             ?@������������������������       �                     7@�       �                   �_@      �?              @������������������������       �                      @�       �                   �b@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   `@���m�?           0{@�       �                    �?�&]�t��?A            �Z@�       �                    �L@      �?0            �S@�       �                   @c@�	j*D�?            �C@������������������������       �                     &@�       �                   8t@h�����?             <@������������������������       �                     :@�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @e@�	j*D�?            �C@�       �       
             �?ҳ�wY;�?             A@�       �                   �l@�+$�jP�?             ;@�       �                    �?�n_Y�K�?             *@������������������������       �                     @�       �                     P@z�G�z�?             $@������������������������       �                     @�       �                    @���Q��?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@������������������������       �                     @������������������������       �                     @�       �                   p`@\-��p�?             =@�       �                   �\@      �?             @������������������������       �                      @������������������������       �                      @�       �       	          pff�?HP�s��?             9@�       �                    �R@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �        	             .@�       �       
             �?"�W1��?�            �t@�       �       
             �?)O���?@             [@������������������������       �                     @�       �                   �f@�7�yHx�?;            @Y@�       �                    �?r�q��?
             2@�       �                    �?�t����?	             1@�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          `ff@��S�ۿ?             .@������������������������       �                     *@�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �l@��a����?1            �T@�       �                    �?      �?             8@�       �                    �?���}<S�?             7@�       �       	             @�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�       �       	          ����?�C��2(�?             &@������������������������       �                     "@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   d@L
�q��?$            �M@�       �                    �?�θ�?            �C@�       �                    �?      �?             0@������������������������       �                     �?������������������������       �                     .@�       �                     N@�LQ�1	�?             7@�       �                    �?؇���X�?             ,@�       �                    �?r�q��?	             (@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �b@ףp=
�?             $@�       �                   @_@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �a@�q�q�?             "@�       �                   �`@z�G�z�?             @�       �       	          Zff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   Pn@      �?             @������������������������       �                     �?�       �                   �y@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   n@�G�z��?             4@�       �                    �?      �?              @�       �                   �e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                     H@r�q��?             (@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�                         �f@P���Q�?�            �k@�       �                    @L@���O�?�            `k@�       �                   @[@���ib#�?t            �e@�       �                    c@�r����?
             .@�       �                    �F@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@������������������������       �        j             d@�       �                   �m@"pc�
�?             F@�       �                   �l@����X�?             5@�       �                    @r�q��?             2@�       �                    _@$�q-�?
             *@������������������������       �                     �?������������������������       �        	             (@�       �       	            �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�                         @a@���}<S�?             7@�                          �M@���Q��?             @                         @d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �        
             2@������������������������       �                     �?�t�b�m(     h�h(h+K ��h-��R�(KMKK��h_�BP       �y@     �@     @Z@     �w@      C@     �s@      ;@      a@      9@     �S@      �?     �F@              ?@      �?      ,@      �?       @               @      �?                      (@      8@      A@      5@      1@      �?       @              @      �?      �?      �?                      �?      4@      "@      $@      �?      @      �?      @                      �?      @              $@       @      @       @      @                       @      @      @      @      �?              �?      @                      @      @      1@      @                      1@       @     �L@              L@       @      �?       @                      �?      &@      f@      @              @      f@      �?     @V@      �?      3@      �?      @              @      �?                      ,@             �Q@      @      V@      @      @      @       @               @      @                      @      @     @T@      �?      @              @      �?               @     �R@      �?      (@      �?      @               @      �?      �?      �?                      �?              "@      �?     �O@              A@      �?      =@      �?      *@      �?                      *@              0@     �P@     @P@      M@      4@       @      @       @      �?              �?       @                      @      L@      .@     �G@       @      *@      @      $@              @      @      @       @      @      �?      �?               @      �?              �?       @                      �?              @      A@       @              �?      A@      �?      @              ;@      �?       @      �?       @                      �?      9@              "@      @      @      @       @      �?       @                      �?       @      @              @       @      �?      �?      �?      �?                      �?      �?              @              "@     �F@      @     �F@      @      0@      �?              @      0@              0@      @               @      =@              7@       @      @               @       @      @              @       @              @             �r@     �`@     �E@      P@     �C@     �C@      ;@      (@              &@      ;@      �?      :@              �?      �?              �?      �?              (@      ;@      (@      6@      @      6@      @       @      @               @       @              @       @      @       @      �?       @                      �?               @              ,@      @                      @      @      9@       @       @               @       @               @      7@       @       @               @       @                      .@     @p@      Q@     �I@     �L@      @              F@     �L@      @      .@       @      .@      �?      �?      �?                      �?      �?      ,@              *@      �?      �?      �?                      �?      �?             �D@      E@      5@      @      5@       @      &@      �?      &@                      �?      $@      �?      "@              �?      �?              �?      �?                      �?      4@     �C@      "@      >@      �?      .@      �?                      .@       @      .@       @      (@       @      $@      �?      �?              �?      �?              �?      "@      �?      @      �?                      @              @               @      @      @      @      �?      �?      �?      �?                      �?      @               @       @      �?              �?       @               @      �?              &@      "@      �?      @      �?       @               @      �?                      @      $@       @       @       @       @                       @       @              j@      &@      j@      $@     �e@       @      *@       @      @       @      @                       @      $@              d@              B@       @      .@      @      .@      @      (@      �?              �?      (@              @       @      @                       @              @      5@       @      @       @      �?       @               @      �?               @              2@                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJѕ:dhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM	hwh(h+K ��h-��R�(KM	��h~�B�9         4                    �?x��X���?=           ��@                          �Q@�9:�l'�?w            @h@������������������������       �                     "@              	          ����?z�G�z�?q             g@                          �s@��a��?K            @^@              
             �?Ц�f*�?C            �[@                          @q@�KM�]�?             3@              	          ����?�X�<ݺ?
             2@	                          �m@      �?             @
                          @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@������������������������       �                     �?                          s@@��,B�?8            �V@������������������������       �        2            �T@                          s@�����H�?             "@������������������������       �                     �?������������������������       �                      @              
             �?���|���?             &@������������������������       �                     @                           �L@      �?              @������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       -                    �M@     ��?&             P@       ,                   �d@��V#�?            �E@       #                   �p@��Q���?             D@                           �n@P���Q�?             4@������������������������       �        
             ,@!       "                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?$       +                    �?      �?             4@%       &                     F@����X�?             ,@������������������������       �                     �?'       *       	          ����?�θ�?             *@(       )                     @      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @.       /                   `l@���N8�?
             5@������������������������       �                     @0       3       	          ����?�IєX�?	             1@1       2                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @5       �                    �?���S��?�           ��@6       k                    @K@�����?�            pz@7       H       
             �?f���oh�?�            �n@8       ;                    �?�0���?-            �T@9       :       	          `ff@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?<       C                   Pr@��a�2��?%             R@=       >                   �h@���#�İ?             �M@������������������������       �                     :@?       @       
             �?�FVQ&�?            �@@������������������������       �                     �?A       B                   �i@      �?             @@������������������������       �                     �?������������������������       �                     ?@D       E                   (s@8�Z$���?             *@������������������������       �                     $@F       G                   `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?I       h                   �g@�G߰K�?^             d@J       _       	          ����?x��-�?\            �c@K       \       	          833�?x�C����?U            �b@L       M                   �k@��<b�ƥ?O            @a@������������������������       �        %            �N@N       Q                   �k@`<)�+�?*            @S@O       P                    b@�q�q�?             @������������������������       �                      @������������������������       �                     �?R       S                   @[@�?�|�?'            �R@������������������������       �                     �?T       [                   `\@ �й���?&            @R@U       V                   �c@�����H�?             "@������������������������       �                     @W       Z                    n@z�G�z�?             @X       Y                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        !             P@]       ^                   �U@z�G�z�?             $@������������������������       �                      @������������������������       �                      @`       g                    �J@�eP*L��?             &@a       b                   �a@      �?              @������������������������       �                      @c       f                   �e@      �?             @d       e                   �l@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @i       j                    �D@      �?              @������������������������       �                     �?������������������������       �                     �?l       �                   �`@v0���1�?r            `f@m       �                   @a@��3E��?7            @W@n                           �?      �?             L@o       |                    �?h+�v:�?             A@p       u       
             �?��<b���?             7@q       r                   `]@      �?             0@������������������������       �                     *@s       t       	          033@�q�q�?             @������������������������       �                     �?������������������������       �                      @v       w                     L@և���X�?             @������������������������       �                      @x       {                   �]@z�G�z�?             @y       z                   @\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @}       ~       	          ����?���!pc�?             &@������������������������       �                      @������������������������       �                     @�       �                    �?���7�?
             6@�       �                    u@��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                     @�       �                    �?�L���?            �B@�       �       	          ����?r�q��?             (@�       �                   `_@�C��2(�?             &@������������������������       �                      @�       �                    `@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �       
             �?`2U0*��?             9@������������������������       �                     6@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?v ��?;            �U@�       �       	          pff�?և���X�?             <@�       �                    �L@     ��?
             0@������������������������       �                     @�       �       	            �?8�Z$���?             *@�       �                    �?�C��2(�?             &@�       �                    �?r�q��?             @�       �                    d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �a@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�       �       
             �?�f7�z�?*             M@�       �                   Pk@�q�q�?             ;@�       �                    �?r�q��?             2@�       �                   �b@�8��8��?             (@�       �                    X@z�G�z�?             @������������������������       �                     @�       �                   b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   0a@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?�n`���?             ?@�       �                    c@����X�?             @������������������������       �                     @������������������������       �                      @�       �                    ]@r�q��?             8@�       �                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    d@�����?             5@�       �                   (p@�}�+r��?             3@������������������������       �        	             (@�       �                     M@؇���X�?             @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?X�EQ]N�?�            �r@�       �                   �`@�'N��?'            �N@�       �                    [@��p\�?            �D@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       
             �?�7��?            �C@������������������������       �                     A@�       �                   @\@���Q��?             @������������������������       �                     @������������������������       �                      @�       �       
             �?�z�G��?             4@������������������������       �                     @�       �                    `@@�0�!��?	             1@������������������������       �                      @�       �                   `d@��S�ۿ?             .@�       �                   �h@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �[@��(\���?�             n@�       �                    �?������?             ;@�       �                     M@�㙢�c�?             7@�       �                    �?������?             .@�       �                    @J@d}h���?
             ,@�       �                   �Z@�8��8��?             (@�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @E@p ��g�?�            �j@�       �                    b@���!pc�?	             &@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                   `U@�q�q�?             @������������������������       �                     �?������������������������       �                      @�                         �e@��'cy�?�            @i@�                         P`@ ���J��?�            `h@�       �       	          ����?      �?.             P@�       �                   8q@      �?             8@������������������������       �                     0@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @�       �       
             �?�(\����?             D@������������������������       �                    �B@�                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �R@��"pK�?R            ``@������������������������       �        P             `@            
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                        �X@և���X�?             @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM	KK��h_�B�       0z@     0@     �b@      G@              "@     �b@     �B@     �\@      @     �Z@      @      1@       @      1@      �?      @      �?      �?      �?      �?                      �?       @              ,@                      �?     �V@      �?     �T@               @      �?              �?       @              @      @              @      @      �?      @               @      �?       @                      �?      A@      >@      =@      ,@      =@      &@      3@      �?      ,@              @      �?      @                      �?      $@      $@      $@      @              �?      $@      @      @      @              @      @              @                      @              @      @      0@      @              �?      0@      �?       @      �?                       @               @     �p@     P|@     �m@     `g@     �e@     �Q@      7@      N@      $@      �?      $@                      �?      *@     �M@       @     �L@              :@       @      ?@      �?              �?      ?@      �?                      ?@      &@       @      $@              �?       @               @      �?             �b@      &@     �b@      $@     �a@      @     �`@      @     �N@             �R@      @       @      �?       @                      �?      R@       @              �?      R@      �?       @      �?      @              @      �?      �?      �?      �?                      �?      @              P@               @       @               @       @              @      @      @      @               @      @      @      @      �?              �?      @                       @      @              �?      �?      �?                      �?     �O@      ]@      1@      S@      ,@      E@      *@      5@      @      2@      �?      .@              *@      �?       @      �?                       @      @      @               @      @      �?      �?      �?      �?                      �?      @               @      @       @                      @      �?      5@      �?      ,@              ,@      �?                      @      @      A@       @      $@      �?      $@               @      �?       @      �?                       @      �?              �?      8@              6@      �?       @      �?                       @      G@      D@      (@      0@      &@      @              @      &@       @      $@      �?      @      �?       @      �?       @                      �?      @              @              �?      �?      �?                      �?      �?      &@      �?                      &@      A@      8@      "@      2@      @      .@      �?      &@      �?      @              @      �?      �?              �?      �?                      @       @      @              @       @      �?              �?       @              @      @      @                      @      9@      @      @       @      @                       @      4@      @      �?       @      �?                       @      3@       @      2@      �?      (@              @      �?      �?      �?              �?      �?              @              �?      �?              �?      �?             �A@     �p@      1@      F@      @      C@      �?      �?              �?      �?               @     �B@              A@       @      @              @       @              ,@      @              @      ,@      @               @      ,@      �?      @      �?              �?      @               @              2@     �k@      @      4@      @      3@      @      &@      @      &@      �?      &@      �?       @               @      �?                      "@       @              �?                       @      @      �?      @                      �?      &@     @i@      @       @      �?      @              @      �?               @      �?              �?       @               @     @h@      @     �g@      @      N@      @      5@              0@      @      @              @      @              �?     �C@             �B@      �?       @      �?                       @      �?     @`@              `@      �?       @      �?                       @      @      @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ1�;hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�5         �       	          ����?b��@�F�?=           ��@       u                    �?(��3�?#           �|@              	          033�dnD��?�            �w@                           �?      �?              @                          �e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @	                          �`@03�Z*!�?�            w@
                           �?������?             �I@                          �_@��2(&�?             F@                          @E@ 7���B�?             ;@������������������������       �                     :@������������������������       �                     �?                          �X@�t����?             1@������������������������       �                     @                           �?�n_Y�K�?
             *@                           @I@�����H�?             "@������������������������       �                     @                          �[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          `Y@؇���X�?             @������������������������       �                     �?������������������������       �                     @       n                   �t@�iʫ{�?�            �s@       E                    �?>a�����?�             s@       <                   �a@\�Uo��?3             S@       7       	          ����?�q�q�?-            �P@       (                   �i@(옄��?             G@        !       
             �?�θ�?             *@������������������������       �                     @"       '                    ^@և���X�?             @#       $                   g@z�G�z�?             @������������������������       �                     �?%       &                   Pa@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @)       *                    �?�q�q�?            �@@������������������������       �                     @+       .                   Xp@�5��?             ;@,       -       
             �?��S�ۿ?             .@������������������������       �                     �?������������������������       �        
             ,@/       6                     M@r�q��?             (@0       1                    �?�C��2(�?             &@������������������������       �                     @2       5                     D@؇���X�?             @3       4                   �a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?8       9                    �?P���Q�?             4@������������������������       �                     1@:       ;                   `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?=       >       
             �?z�G�z�?             $@������������������������       �                     @?       D                   �d@����X�?             @@       A                   �b@r�q��?             @������������������������       �                     @B       C                    �G@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?F       Y                    �?ج��w�?�            �l@G       N                    �?�<ݚ�?             B@H       M                   �`@      �?              @I       J                    @L@���Q��?             @������������������������       �                      @K       L       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @O       V                   �q@ �Cc}�?             <@P       Q       	          pff�?$�q-�?             :@������������������������       �                     3@R       S                   �_@����X�?             @������������������������       �                     @T       U       	          ����?      �?             @������������������������       �                      @������������������������       �                      @W       X                   s@      �?              @������������������������       �                     �?������������������������       �                     �?Z       k                    �?h�a��?{            @h@[       h                    @`k�����?k             e@\       g                    �?�O4R���?c            �c@]       ^                   Pn@��<b�ƥ?U            @a@������������������������       �        2             U@_       b       
             �?�X�<ݺ?#             K@`       a                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?c       f                   @[@���J��?!            �I@d       e                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �H@������������������������       �                     5@i       j       
             �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @l       m       
             �?���B���?             :@������������������������       �                     @������������������������       �                     5@o       t                    �M@      �?             (@p       s                    �?      �?              @q       r       
             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @v       y                    [@U7W1�?/            �T@w       x       	             �r�q��?             @������������������������       �                     �?������������������������       �                     @z       �       
             �?6��f�?,            @S@{       �                   �b@$�q-�?             J@|       �                    �?`2U0*��?             I@}       �                    �K@�FVQ&�?            �@@~       �                   �l@�q�q�?             @       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     ;@������������������������       �        	             1@������������������������       �                      @�       �                    I@�q�����?             9@������������������������       �                     @�       �                    �H@p�ݯ��?	             3@������������������������       �                     @�       �                   �h@؇���X�?             ,@�       �                   �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     $@�       �       	          ���@�t����?           �|@�       �                   �b@ kGZ=��?�            0v@�       �                    �?�LQ�1	�?�            @q@�       �                    �?�G��l��?             E@�       �                    `@�\��N��?             C@�       �                   �\@�E��ӭ�?             2@�       �                    �L@����X�?             @�       �                   Pp@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     &@�       �                    @K@��Q��?             4@�       �                   n@��
ц��?	             *@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?|�űN�?�            @m@�       �                   `S@r�q��?#             N@������������������������       �                      @�       �       
             �?\-��p�?"             M@�       �                    �?��S�ۿ?            �F@�       �                   �k@z�G�z�?             $@������������������������       �                     @�       �       
             �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �a@��?^�k�?            �A@������������������������       �                     <@�       �       	             �?؇���X�?             @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �a@�n_Y�K�?             *@������������������������       �                      @������������������������       �                     @�       �                    �R@XB���?o            �e@�       �                   j@������?m            �e@�       �                    �?$�q-�?,            @P@�       �                    �M@     ��?             @@�       �       	          ����?�C��2(�?             6@�       �                   @Y@�r����?             .@������������������������       �                     �?�       �                   �c@@4և���?             ,@������������������������       �                     "@�       �                   �f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �d@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                    �@@������������������������       �        A            �Z@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @L@v�_���?3            �S@�       �       	          ����?��k=.��?             �G@�       �                    �?և���X�?	             ,@������������������������       �                      @�       �                    �?      �?             (@������������������������       �                     @�       �                    �?؇���X�?             @������������������������       �                     @�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `T@�C��2(�?            �@@������������������������       �                     �?�       �                   �e@      �?             @@������������������������       �                     9@�       �       	             �?����X�?             @������������������������       �                     @�       �                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?     ��?             @@�       �                    �?j���� �?	             1@������������������������       �                     $@������������������������       �                     @�       �                    @O@������?
             .@�       �                   `b@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                   pc@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?�]��?7            �Y@�       �                   �Z@ ���J��?)            �S@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        '            �R@�       �                   �c@HP�s��?             9@������������������������       �                     6@�       �       	          033@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       `x@     ��@     �r@     @d@     Pq@      Y@      �?      @      �?      @              @      �?                      @     @q@     @W@      (@     �C@      @      C@      �?      :@              :@      �?              @      (@              @      @       @      �?       @              @      �?      @      �?                      @      @              @      �?              �?      @             �p@      K@      p@      H@      G@      >@      F@      6@      9@      5@      @      $@              @      @      @      �?      @              �?      �?      @      �?                      @       @              6@      &@      @              0@      &@      ,@      �?              �?      ,@               @      $@      �?      $@              @      �?      @      �?      @      �?                      @              @      �?              3@      �?      1@               @      �?       @                      �?       @       @              @       @      @      �?      @              @      �?       @               @      �?              �?             �j@      2@      <@       @      @      @      @       @       @              �?       @               @      �?                      @      9@      @      8@       @      3@              @       @      @               @       @               @       @              �?      �?              �?      �?              g@      $@     `d@      @     �c@      @     �`@      @      U@             �I@      @      �?       @               @      �?              I@      �?      �?      �?              �?      �?             �H@              5@              @       @               @      @              5@      @              @      5@              @      @      @       @      @      �?              �?      @                      �?              @      5@      O@      @      �?              �?      @              0@     �N@      @      H@       @      H@       @      ?@       @      @       @      �?       @                      �?              @              ;@              1@       @              (@      *@              @      (@      @              @      (@       @       @       @       @                       @      $@              W@     �v@      V@     �p@      B@      n@      4@      6@      4@      2@      *@      @       @      @       @      �?              �?       @                      @      &@              @      *@      @      @      @               @      @              @       @                      @              @      0@     @k@      $@      I@       @               @      I@      @      E@       @       @              @       @      @       @                      @      �?      A@              <@      �?      @      �?      �?      �?                      �?              @      @       @               @      @              @      e@      @     �d@      @      N@      @      ;@       @      4@       @      *@      �?              �?      *@              "@      �?      @      �?                      @              @      @      @              @      @                     �@@             �Z@      �?      �?      �?                      �?      J@      ;@      C@      "@       @      @       @              @      @              @      @      �?      @              �?      �?              �?      �?              >@      @              �?      >@       @      9@              @       @      @              �?       @      �?                       @      ,@      2@      $@      @      $@                      @      @      &@      �?       @               @      �?              @      @      @                      @      @     �X@       @      S@       @      �?       @                      �?             �R@       @      7@              6@       @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ'�ShG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�9         �                    �?<qn�h��?=           ��@       -                    _@ x�Y��?`           �@                           �?�2�IQ�?;            �V@       	       
             �?      �?)             P@                           �?��Y��]�?            �D@������������������������       �                     >@              
             �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@
                          �^@8����?             7@                           \@X�<ݚ�?             "@������������������������       �                     @                           �J@z�G�z�?             @������������������������       �                     �?������������������������       �                     @              	          `ff�?؇���X�?	             ,@              	             �?���Q��?             @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     "@       ,                     R@
j*D>�?             :@       #       	          ����?      �?             6@              	             ���<ݚ�?             "@������������������������       �                     @       "                   �^@�q�q�?             @       !       
             �?      �?             @                           \@�q�q�?             @������������������������       �                     �?                            @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @$       %                    @J@�	j*D�?	             *@������������������������       �                      @&       '                    �?"pc�
�?             &@������������������������       �                     @(       )                    �?�q�q�?             @������������������������       �                      @*       +                   @c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @.       �       	          ���@�1f����?%           �|@/       l                    �J@"�R�}q�?           �{@0       I                   �]@J�:�Ȣ�?�            �o@1       F                    ]@�BbΊ�?*             M@2       E                   @f@��x_F-�?$            �I@3       :                     D@��[�p�?             �G@4       5                    @A@      �?             $@������������������������       �                     @6       7                    @C@����X�?             @������������������������       �                     @8       9                   �a@      �?             @������������������������       �                      @������������������������       �                      @;       @                   Hp@$G$n��?            �B@<       =       
             �?`Jj��?             ?@������������������������       �                     �?>       ?                    f@(;L]n�?             >@������������������������       �                     =@������������������������       �                     �?A       D                    �?      �?             @B       C                   0`@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @G       H                   b@����X�?             @������������������������       �                     @������������������������       �                      @J       _       
             �?�q��/��?            �h@K       V                   ``@��S���?            �F@L       U                    �?8^s]e�?             =@M       N                   �f@�θ�?             :@������������������������       �                     �?O       T                    �?z�G�z�?             9@P       S                   �q@�q�q�?             (@Q       R                    �I@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        	             *@������������������������       �                     @W       X                    �?      �?
             0@������������������������       �                     �?Y       \                   �e@z�G�z�?	             .@Z       [                    �E@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@]       ^                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @`       k                    �? Gn���?c            �b@a       b                    �?ȵHPS!�?             :@������������������������       �                      @c       j                   Hp@r�q��?             2@d       i                   �n@      �?	             (@e       h       	             �?"pc�
�?             &@f       g                   @b@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        O            @_@m       �                    c@�_;"�?t            `g@n       �       
             �?r�u���?e            �d@o       p       	          833�?X�<ݚ�?'            �O@������������������������       �        
             2@q       �                   �r@F�����?            �F@r       u       	          ����?��%��?            �B@s       t                    �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?v       {                    �?�5��?             ;@w       x       	          033�?���Q��?             $@������������������������       �                      @y       z                    �?      �?              @������������������������       �                     @������������������������       �                      @|       }                   �h@�t����?             1@������������������������       �                      @~                          �b@z�G�z�?
             .@������������������������       �                     "@�       �                    �?      �?             @�       �                   `c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �?ȵHPS!�?>             Z@�       �                    �?���|���?             6@�       �       	            �?D�n�3�?             3@�       �                   �b@d}h���?
             ,@������������������������       �                      @�       �                   �c@      �?             @������������������������       �                      @�       �                    �?      �?             @�       �                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?������?1            �T@�       �                    @L@�X�<ݺ?)             R@������������������������       �                     ?@�       �                   p@������?            �D@������������������������       �                     7@�       �                    �?�<ݚ�?
             2@�       �       	          ����?X�<ݚ�?             "@�       �                    @M@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �                     $@�       �                   �c@�z�G��?             4@�       �                    �?      �?             (@������������������������       �                     @�       �                    @N@�q�q�?             "@�       �                    X@���Q��?             @������������������������       �                      @�       �                   `n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �]@�r����?             .@������������������������       �                      @������������������������       �                     *@�       �                    �?�T�p �?�            @w@�       �       
             �?H�z�G�?             D@�       �                    �?     ��?             @@�       �       	          ����?և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �`@z�G�z�?             9@�       �                   u@X�Cc�?             ,@�       �                   �k@z�G�z�?             $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                      @�       �                    �?\�>���?�            �t@�       �                    Z@0�v���?�            `p@�       �       	             @�eP*L��?             &@�       �                   0a@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �R@`�ҕ�ļ?�            `o@�       �                   pa@�>��(+�?�             o@�       �                   �\@0�z��?�?J             _@�       �                    @L@ >�֕�?            �A@������������������������       �                     1@�       �                    �?�����H�?             2@������������������������       �        	             &@�       �       
             �?����X�?             @�       �                   �^@r�q��?             @������������������������       �                     @�       �                   �Y@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �        1            @V@�       �                   �b@����y7�?J            @_@�       �       
             �?@4և���?D             \@�       �                     E@ }�Я��?7            @V@�       �                    `@      �?             @�       �                    �C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        4            @U@�       �                   `j@8����?             7@�       �                    c@ףp=
�?             $@������������������������       �                      @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?��
ц��?             *@������������������������       �                     @������������������������       �                     @�       �                    n@�	j*D�?             *@������������������������       �                      @�       �                   �b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �h@��R[s�?*            �Q@�       �                   @e@(;L]n�?             >@������������������������       �                     =@������������������������       �                     �?�             
             �?H�z�G�?             D@�                         �b@V�a�� �?             =@�       �                   �\@H%u��?             9@������������������������       �                     �?�                          �s@�8��8��?             8@�       �                    @N@���7�?             6@������������������������       �                     (@�       �                   �`@ףp=
�?             $@������������������������       �                     @�       �                     P@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �K@      �?              @������������������������       �                     �?������������������������       �                     �?            	          033@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KMKK��h_�Bp       z@     P@     �v@      g@      3@     �Q@       @      L@      �?      D@              >@      �?      $@      �?                      $@      @      0@      @      @      @              �?      @      �?                      @       @      (@       @      @      �?      @      �?                      @      �?                      "@      &@      .@      &@      &@       @      @              @       @      @       @       @      �?       @              �?      �?      �?              �?      �?              �?                       @      "@      @               @      "@       @      @              @       @       @               @       @               @       @                      @     pu@     @\@     Pu@      Y@     �j@     �C@     �E@      .@     �D@      $@     �B@      $@      @      @      @               @      @              @       @       @       @                       @      @@      @      =@       @              �?      =@      �?      =@                      �?      @      @      @       @      @                       @              �?      @               @      @              @       @             �e@      8@      8@      5@      4@      "@      4@      @              �?      4@      @      @      @      �?      @              @      �?              @              *@                      @      @      (@      �?              @      (@      �?      &@      �?                      &@       @      �?              �?       @             �b@      @      7@      @       @              .@      @      "@      @      "@       @      "@      �?      "@                      �?              �?              �?      @             @_@             �_@     �N@      ^@     �G@      <@     �A@              2@      <@      1@      4@      1@      "@      �?      "@                      �?      &@      0@      @      @               @      @       @      @                       @      @      (@       @              @      (@              "@      @      @      �?      @      �?                      @       @               @              W@      (@      ,@       @      &@       @      &@      @       @              @      @               @      @      �?       @      �?       @                      �?      �?                      @      @             �S@      @      Q@      @      ?@             �B@      @      7@              ,@      @      @      @      @      @              @      @               @              "@              $@              @      ,@      @      @              @      @      @       @      @               @       @      �?       @                      �?      @                       @       @      *@       @                      *@     �K@     �s@      1@      7@      "@      7@      @      @      @                      @      @      4@      @      "@       @       @              @       @      @       @                      @      @      �?      @                      �?              &@       @              C@     `r@      4@     @n@      @      @      �?      @              @      �?              @              .@     �m@      ,@     `m@       @     �^@       @     �@@              1@       @      0@              &@       @      @      �?      @              @      �?       @               @      �?              �?                     @V@      (@     @\@       @      Z@      �?      V@      �?      @      �?      �?              �?      �?                       @             @U@      @      0@      �?      "@               @      �?      �?              �?      �?              @      @      @                      @      @      "@               @      @      �?      @                      �?      �?      �?      �?                      �?      2@      J@      �?      =@              =@      �?              1@      7@      @      7@      @      6@      �?               @      6@      �?      5@              (@      �?      "@              @      �?       @      �?                       @      �?      �?              �?      �?              @      �?      @                      �?      &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJŮ�dhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM	hwh(h+K ��h-��R�(KM	��h~�B�9         �                    �?��J�0�?Q           ��@       ]       
             �?|z U���?Z           ��@       X                    �?������?�            �w@                          �Z@\-��p�?�            Pp@              
             �?      �?              @������������������������       �                      @                           �?�q�q�?             @������������������������       �                     @	       
                    �D@�q�q�?             @������������������������       �                     �?                          �o@      �?              @������������������������       �                     �?������������������������       �                     �?       I                   �b@��FƘ��?�            �o@       H                     P@���}<S�?�            �l@                           �?����#��?�             i@                           �?�LQ�1	�?             7@                          �`@�X����?             6@                          �_@����X�?             @������������������������       �                     �?                           �I@r�q��?             @������������������������       �                     �?������������������������       �                     @                          �`@�r����?	             .@              	             �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?       C                    �O@���M�?t            @f@       .                   `_@�}�+r��?p            `e@        '       	             @@��8��?B             X@!       &                   `P@�Fǌ��?7            �S@"       #                    @O@(;L]n�?             >@������������������������       �                     ;@$       %                   �Y@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        #            �H@(       )       
             �?�IєX�?             1@������������������������       �                      @*       -                   ``@��S�ۿ?
             .@+       ,                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@/       4                    \@���Lͩ�?.            �R@0       1       	             �?���Q��?             $@������������������������       �                     @2       3                   �a@և���X�?             @������������������������       �                     @������������������������       �                     @5       <                   `h@P�2E��?(            @P@6       9                    @G@"pc�
�?             &@7       8                    `@�q�q�?             @������������������������       �                     �?������������������������       �                      @:       ;                   `g@      �?              @������������������������       �                     @������������������������       �                     �?=       B                    �H@@3����?!             K@>       ?                   �p@�C��2(�?             &@������������������������       �                      @@       A                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �E@D       G       	             �?և���X�?             @E       F                    j@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     =@J       M                   Po@\X��t�?             7@K       L                   pd@�q�q�?             "@������������������������       �                     @������������������������       �                     @N       Q                    �?����X�?
             ,@O       P       	             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @R       S       	          ����?���Q��?             @������������������������       �                      @T       W                    �?�q�q�?             @U       V                   0c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?Y       Z                   �c@ 4^��?O            �]@������������������������       �        ?             X@[       \                   �r@�nkK�?             7@������������������������       �                     6@������������������������       �                     �?^       �                    �?D����?`            �b@_       z                    �L@d��0u��?L             ^@`       c                   @E@��W��?/            @R@a       b                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @d       e                    �?��hJ,�?,             Q@������������������������       �                     5@f       s       	          433�?��[�p�?             �G@g       r                    �?      �?             D@h       q                   �b@�חF�P�?             ?@i       j                   �c@ܷ��?��?             =@������������������������       �                     1@k       l                   @i@      �?	             (@������������������������       �                      @m       n                    �?ףp=
�?             $@������������������������       �                     @o       p                    ]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     "@t       y                    �?����X�?             @u       v                   0e@r�q��?             @������������������������       �                     @w       x                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?{       �                   �r@Z�K�D��?            �G@|       �                   �e@�s��:��?             C@}       �       	          ����?���Q��?            �A@~       �                    �?b�2�tk�?             2@       �                   �l@      �?	             (@�       �       	          ����?�q�q�?             "@�       �                    �?���Q��?             @�       �                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �[@r�q��?             @�       �                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    c@@�0�!��?             1@������������������������       �                     ,@������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �       	          ����?ܷ��?��?             =@�       �                   ``@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     6@�       �                   �_@Z�EΡ-�?�            Px@�       �                    �?���j��?             G@�       �                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                   �e@4?,R��?             B@�       �                   �c@�C��2(�?            �@@�       �       
             �?XB���?             =@������������������������       �                     :@�       �       	          ����?�q�q�?             @������������������������       �                     �?�       �                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �F@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @N@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   `@�ӝ��?�            pu@�       �       
             �?�ݜ����?(            �M@�       �                     P@ףp=
�?             >@������������������������       �                     8@�       �                    `Q@      �?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �p@\-��p�?             =@������������������������       �                     7@�       �       	          hff�?�q�q�?             @�       �                   �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�             	          ���@�������?�            �q@�       �       
             �?�㙢�c�?�            @q@�       �                   `a@�q�����?/            �R@�       �                    �B@�LQ�1	�?             G@������������������������       �                     @�       �       	          ����?�^�����?            �E@�       �                    �?�eP*L��?             &@�       �                    �J@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �g@      �?             @@�       �                   �b@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�>4և��?             <@�       �                   @q@�q�q�?             (@�       �       	          033�?�����H�?             "@�       �       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          ����?      �?             0@�       �                    �K@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             (@�       �       	          ����?V�a�� �?             =@�       �                     Q@�KM�]�?             3@�       �                    @�X�<ݺ?
             2@�       �                    b@@4և���?             ,@������������������������       �                      @�       �                   pl@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �c@���Q��?             $@�       �       	          ����?�q�q�?             @������������������������       �                      @�       �                    �N@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   �l@�����?}             i@������������������������       �        ;            �X@�                         �g@l��\��?B            �Y@�                         �d@D���ͫ�?A            @Y@�       �                   �n@\-��p�?$             M@�       �       	          ����?��
ц��?             *@�       �                    �?�q�q�?             "@������������������������       �                      @�       �                    �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?`Ӹ����?            �F@������������������������       �                     2@�       �                    _@�>����?             ;@�       �                    �K@؇���X�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?                          �O@P���Q�?             4@������������������������       �        
             2@                        Pb@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �E@������������������������       �                     �?                        �f@      �?              @������������������������       �                     @������������������������       �                     �?�t�b�     h�h(h+K ��h-��R�(KM	KK��h_�B�        x@     ��@      ]@     �y@     �B@     pu@      B@      l@      @       @       @              @       @      @              �?       @              �?      �?      �?      �?                      �?      >@     �k@      4@     @j@      4@     �f@       @      .@      @      .@      @       @              �?      @      �?              �?      @               @      *@       @      @       @                      @               @      �?              (@     �d@      "@     @d@       @     �W@      �?     �S@      �?      =@              ;@      �?       @               @      �?                     �H@      �?      0@               @      �?      ,@      �?       @               @      �?                      (@      @      Q@      @      @              @      @      @      @                      @      @      O@       @      "@      �?       @      �?                       @      �?      @              @      �?              �?     �J@      �?      $@               @      �?       @      �?                       @             �E@      @      @      @      �?              �?      @                      @              =@      $@      *@      @      @      @                      @      @      $@      �?       @      �?                       @      @       @       @              �?       @      �?      �?              �?      �?                      �?      �?     �]@              X@      �?      6@              6@      �?             �S@     �Q@      S@      F@     �M@      ,@      �?      @      �?                      @      M@      $@      5@             �B@      $@     �A@      @      :@      @      :@      @      1@              "@      @               @      "@      �?      @              @      �?              �?      @                       @      "@               @      @      �?      @              @      �?      �?      �?                      �?      �?              1@      >@      1@      5@      ,@      5@      &@      @      @      @      @      @       @      @       @      �?       @                      �?               @      @                      @      @      �?       @      �?       @                      �?      @              @      ,@              ,@      @              @                      "@      @      :@      @      @              @      @                      6@     �p@     �]@      *@     �@@       @       @       @                       @      @      ?@      @      >@      �?      <@              :@      �?       @              �?      �?      �?              �?      �?               @       @      �?              �?       @              �?      �?      �?      �?                      �?       @      �?       @                      �?     p@     �U@      <@      ?@      @      ;@              8@      @      @       @              �?      @              @      �?              9@      @      7@               @      @       @       @       @                       @               @     �l@     �K@     �l@      H@      B@     �C@      >@      0@              @      >@      *@      @      @      @      �?      @                      �?              @      8@       @      �?      @      �?                      @      7@      @       @      @       @      �?      @      �?              �?      @              @                      @      .@      �?      @      �?      @                      �?      (@              @      7@       @      1@      �?      1@      �?      *@               @      �?      @              @      �?                      @      �?              @      @      @       @       @               @       @       @                       @              @      h@      "@     �X@             @W@      "@     @W@       @      I@       @      @      @      @      @               @      @      @      @                      @      @             �E@       @      2@              9@       @      @      �?      @              �?      �?              �?      �?              3@      �?      2@              �?      �?      �?                      �?     �E@                      �?      �?      @              @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ&��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B�4         �                    �?�lb���?L           ��@                          `X@�%�a�u�?_           ��@������������������������       �                     @       K       
             �?q�H5�?[           ��@                           �?�����?�            �i@                           �O@� �	��?!             I@                           �?      �?             F@                          �a@ҳ�wY;�?             A@	       
                   �Q@�+$�jP�?             ;@������������������������       �                     �?                          �]@8�Z$���?             :@������������������������       �                     (@                          l@����X�?             ,@������������������������       �                     @                           e@      �?              @                           �?�q�q�?             @������������������������       �                      @                           �K@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     $@������������������������       �                     @               
             �?Tݭg_�?c            �c@                          e@      �?             0@                           �?���!pc�?             &@������������������������       �                     @                           `Q@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @!       J                   @f@R���Q�?X            �a@"       -       	          ����?d/�@7�?V             a@#       $                    �?h�����?%             L@������������������������       �                    �D@%       ,                    j@�r����?             .@&       +                   �a@����X�?             @'       (                    @H@�q�q�?             @������������������������       �                     �?)       *                   `X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @.       I                    �Q@|��"J�?1            @T@/       <       	          ����?��t���?0            �S@0       1                    X@�\��N��?             3@������������������������       �                     @2       9                    �?�q�q�?	             .@3       8                    �?�����H�?             "@4       5       	          ����?�q�q�?             @������������������������       �                     �?6       7                   Po@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @:       ;                     @�q�q�?             @������������������������       �                     @������������������������       �                      @=       F                   pr@��S�ۿ?$             N@>       ?                    d@�8���?"             M@������������������������       �                     H@@       E                    �?�z�G��?             $@A       B                    ]@և���X�?             @������������������������       �                      @C       D                   xp@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @G       H                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @L       m                    �L@�����b�?�            @v@M       d                    �?��!���?�             q@N       S                    P@4�2%ޑ�?*            �Q@O       P                    �?ףp=
�?             $@������������������������       �                     @Q       R                   `[@�q�q�?             @������������������������       �                     �?������������������������       �                      @T       W                    @D@�?�P�a�?#             N@U       V                   @b@�z�G��?             $@������������������������       �                     @������������������������       �                     @X       _                   �d@HP�s��?             I@Y       Z                   �b@�(\����?             D@������������������������       �                     @@[       ^                    �G@      �?              @\       ]                    �E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @`       a                    �?�z�G��?             $@������������������������       �                     �?b       c                   `k@�q�q�?             "@������������������������       �                     @������������������������       �                     @e       l       	             @0���{�?y            �i@f       i                    @L@���9�,�?x             i@g       h                   0h@��O{��?u            �h@������������������������       �        t            �h@������������������������       �                     �?j       k                   Hp@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @n       u                    @M@#z�i��?4            �T@o       t       	          ����?�q�q�?             8@p       s                    �?�q�q�?             (@q       r                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@v       �                     R@V�a�� �?(             M@w       �       	          ���@�iʫ{�?%            �J@x                          �c@H%u��?$             I@y       ~                    �M@Pa�	�?            �@@z       {                   `c@؇���X�?             @������������������������       �                     @|       }                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     :@�       �                    �M@�t����?             1@�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �r@d}h���?	             ,@�       �                    �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                   @^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �a@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       
             �?d�|D���?�            �u@�       �                    �? i���t�?�            `r@�       �                   �b@�D�����?�            @k@�       �                    �M@�qM�R��?�             i@�       �                   �Z@ ����?Z            ``@�       �       	          ����?      �?             @������������������������       �                     �?�       �                    �D@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    @K@ d��u�?U            @_@�       �                    `@ >�֕�?2            �Q@������������������������       �        $             J@�       �                    �?�<ݚ�?             2@�       �                    �F@����X�?             ,@������������������������       �                     @�       �                   @b@և���X�?             @�       �       	             �?�q�q�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    `@"pc�
�?#            �K@�       �       	          ����?�E��ӭ�?             B@�       �                   �]@     ��?             0@�       �                   �[@���|���?             &@�       �                    d@և���X�?             @�       �       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   `_@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �                     3@�       �                   ``@`����֜?-            �Q@�       �                   �_@ �q�q�?             8@������������������������       �                     0@�       �                    �?      �?              @�       �                   `]@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     G@�       �                    �?��.k���?	             1@������������������������       �                     @�       �                    �?z�G�z�?             $@������������������������       �                     @�       �                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    @N@p�|�i�?4             S@������������������������       �        "             J@�       �                   �`@      �?             8@�       �                   �Y@P���Q�?             4@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@�       �                   `^@      �?             @������������������������       �                     �?�       �                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          pff�?և���X�?)             L@�       �                     O@j���� �?             A@�       �                    �?��X��?             <@�       �                    h@      �?             2@������������������������       �                     @�       �                    @J@X�Cc�?             ,@�       �                   `m@      �?              @������������������������       �                     �?�       �                   0a@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?"pc�
�?             6@�       �                    �?�KM�]�?             3@�       �                    c@"pc�
�?	             &@�       �                   �`@ףp=
�?             $@�       �                    �M@z�G�z�?             @������������������������       �                      @�       �                    �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B        z@     @@     �v@     �i@              @     �v@     �h@     �L@     �b@      <@      6@      6@      6@      6@      (@      6@      @              �?      6@      @      (@              $@      @      @              @      @      @       @       @               @       @       @                       @               @              @              $@      @              =@     �_@       @       @      @       @              @      @      �?      @                      �?      @              5@     �]@      2@     �]@       @      K@             �D@       @      *@       @      @       @      �?      �?              �?      �?      �?                      �?              @               @      0@     @P@      ,@     @P@      $@      "@              @      $@      @       @      �?       @      �?      �?              �?      �?      �?                      �?      @               @      @              @       @              @      L@      @     �K@              H@      @      @      @      @               @      @       @      @                       @              @      �?      �?              �?      �?               @              @             0s@     �H@     �o@      5@      K@      0@      �?      "@              @      �?       @      �?                       @     �J@      @      @      @      @                      @      G@      @     �C@      �?      @@              @      �?      �?      �?      �?                      �?      @              @      @      �?              @      @              @      @             �h@      @     �h@       @     �h@      �?     �h@                      �?       @      �?       @                      �?              @      K@      <@       @      0@       @      @      �?      @              @      �?              @                      (@      G@      (@      F@      "@      F@      @      @@      �?      @      �?      @               @      �?              �?       @              :@              (@      @      �?       @      �?                       @      &@      @      $@      �?      $@                      �?      �?       @      �?                       @              @       @      @       @                      @      K@     �r@      >@     �p@      ;@     �g@      2@     �f@      1@     �\@      @      @              �?      @       @               @      @              ,@     �[@      @     �P@              J@      @      ,@      @      $@              @      @      @      @       @      @              �?       @               @      �?                      �?              @      $@     �F@      $@      :@      "@      @      @      @      @      @      @      �?              �?      @                       @              @      @              �?      3@              3@      �?                      3@      �?     @Q@      �?      7@              0@      �?      @      �?      @              @      �?                       @              G@      "@       @      @               @       @              @       @      @       @                      @      @     @R@              J@      @      5@      �?      3@      �?      @              @      �?                      0@       @       @              �?       @      �?       @                      �?      8@      @@      4@      ,@      3@      "@      "@      "@              @      "@      @      @      @      �?               @      @       @                      @      @              $@              �?      @              @      �?              @      2@       @      1@       @      "@      �?      "@      �?      @               @      �?       @      �?                       @              @      �?                       @       @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJb�pMhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�5         �       
             �?��.k���?G           ��@                           e@�fC���?A           `@                           �F@��.N"Ҭ?Q            @a@                          �Q@r�q��?             @������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?	                           �?`���i��?L            �`@
                          �a@@��!�Q�?9            @Z@������������������������       �        /            �V@                           �J@@4և���?
             ,@                            J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@                           @O@�>����?             ;@                          @e@�nkK�?             7@������������������������       �                     5@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?              
             �?      �?             @������������������������       �                      @                          �a@      �?              @������������������������       �                     �?������������������������       �                     �?       �       	          ���@�:���?�            �v@       X                    �?6�N���?�            �r@       S                    �?��:#�|�?            �g@       ,                    �?v���a�?d            @b@        %                    �?�LQ�1	�?             7@!       "                    �?      �?             @������������������������       �                      @#       $                   �n@      �?              @������������������������       �                     �?������������������������       �                     �?&       '                   �_@�d�����?             3@������������������������       �                     @(       )                   pl@�q�q�?	             .@������������������������       �                     @*       +       	          ����?r�q��?             (@������������������������       �                      @������������������������       �                     $@-       @                   �`@����X��?S            �^@.       /                    @H@ >�֕�?1            �Q@������������������������       �                     :@0       ?       	             �?�C��2(�?              F@1       >                    a@\-��p�?             =@2       7                   `_@z�G�z�?             4@3       6       	          ����?@4և���?
             ,@4       5       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@8       =                   Pt@      �?             @9       :                    �H@      �?             @������������������������       �                      @;       <                   0j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     .@A       B                   `h@r�����?"            �J@������������������������       �                     @C       R                    `R@�:pΈ��?              I@D       E                    �?dP-���?            �G@������������������������       �                     &@F       I                   �`@�����H�?             B@G       H                    �I@�q�q�?             @������������������������       �                     @������������������������       �                      @J       Q                    c@��S�ۿ?             >@K       P                    �?XB���?             =@L       M                    @K@�nkK�?             7@������������������������       �                     2@N       O                   �a@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @T       W                    �G@�Ń��̧?             E@U       V                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     D@Y       �                    �?�eP*L��?G            �[@Z       _       
             �?L�uϪ�?>            �X@[       ^                    @I@@4և���?             ,@\       ]                    �G@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@`       s                    @K@��6���?7             U@a       b                   �a@�<ݚ�?             B@������������������������       �                     @c       d                    �F@      �?             @@������������������������       �                     &@e       f                    �?��s����?             5@������������������������       �                      @g       n                    �H@�	j*D�?
             *@h       m                    �?      �?             @i       l                    �?�q�q�?             @j       k                     H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?o       r       	          ����?�����H�?             "@p       q                   �j@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @t       }                    �?      �?             H@u       |                    �?���|���?	             &@v       w                   `X@�z�G��?             $@������������������������       �                      @x       {                   �b@      �?              @y       z                    @L@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?~       �                   o@V������?            �B@       �                    �?ҳ�wY;�?
             1@������������������������       �                     @�       �                    `P@      �?             (@�       �                   �b@      �?              @������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@�       �                    �?�8��8��?	             (@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �       	          `ff@Pa�	�?*            �P@�       �                    �? ������?(            �O@������������������������       �                     $@�       �                    �?�O4R���?             �J@������������������������       �                    �C@�       �                     K@@4և���?             ,@�       �       	             @r�q��?             @�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?������?            z@�       �                    �?���)�?T             a@�       �                   �Z@�I� �?8             W@������������������������       �                     @�       �                   �a@���?6            @V@�       �                    U@�ݜ�?            �C@������������������������       �                     �?�       �                   @E@�KM�]�?             C@������������������������       �                     @������������������������       �                     A@�       �                    �?� �	��?             I@�       �                   `\@F�����?            �F@������������������������       �                     @�       �                    �?�(�Tw��?            �C@�       �                    s@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�       �                   @b@��X��?             <@������������������������       �                     @�       �                    �?�+e�X�?             9@�       �                   @f@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   pf@���y4F�?
             3@������������������������       �        	             .@������������������������       �                     @������������������������       �                     @�       �                   (p@�zv�X�?             F@�       �                    @N@�������?             >@�       �                    �?��Q��?             4@�       �                    �?��
ц��?	             *@������������������������       �                     @�       �                    V@���Q��?             $@�       �                    �?���Q��?             @�       �                   �X@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �I@z�G�z�?             @�       �                   pj@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     $@�       �                   �p@����X�?             ,@������������������������       �                     @�       �                    �?X�<ݚ�?             "@������������������������       �                     @�       �                    @J@�q�q�?             @�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          ���@ >�֕�?�            �q@�       �                    @L@`2U0*��?�            0q@�       �       	             �?@p�<��?�             k@������������������������       �        z            �h@�       �                    �?P���Q�?             4@�       �                   �g@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@�       �                    �?�:�B��?&            �M@�       �                   Hs@�C��2(�?             6@�       �                   `b@���N8�?             5@������������������������       �                     3@�       �                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �       	          `ff�?���@��?            �B@�       �                   `a@b�h�d.�?            �A@������������������������       �        	             1@�       �                    �Q@�q�q�?             2@�       �                     P@      �?             0@�       �                    �?���Q��?             $@�       �                    �?      �?              @������������������������       �                     @�       �                   @e@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP        {@     `~@     @V@     �y@      @     �`@      �?      @              @      �?      �?      �?                      �?      @      `@      �?      Z@             �V@      �?      *@      �?      �?              �?      �?                      (@       @      9@      �?      6@              5@      �?      �?              �?      �?              �?      @               @      �?      �?              �?      �?             @U@     pq@     �T@     �j@      7@     �d@      6@      _@       @      .@      @      �?       @              �?      �?      �?                      �?      @      ,@              @      @      $@      @               @      $@       @                      $@      ,@     @[@      @     �P@              :@      @      D@      @      9@      @      0@      �?      *@      �?       @               @      �?                      &@      @      @      @      �?       @              �?      �?      �?                      �?               @              "@              .@      $@     �E@      @              @     �E@      @     �E@              &@      @      @@       @      @              @       @               @      <@      �?      <@      �?      6@              2@      �?      @      �?                      @              @      �?              @              �?     �D@      �?      �?              �?      �?                      D@      N@      I@     �M@     �C@      *@      �?       @      �?       @                      �?      &@              G@      C@      <@       @              @      <@      @      &@              1@      @       @              "@      @      �?      @      �?       @      �?      �?      �?                      �?              �?              �?       @      �?      @      �?      @                      �?      @              2@      >@      @      @      @      @               @      @      �?      @      �?              �?      @              @                      �?      &@      :@      &@      @      @              @      @      @       @      @              �?       @               @      �?                      @              4@      �?      &@      �?      �?              �?      �?                      $@       @      P@      �?      O@              $@      �?      J@             �C@      �?      *@      �?      @      �?      @      �?                      @               @               @      �?       @      �?                       @     pu@     @R@     �S@     �L@      O@      >@              @      O@      ;@      A@      @              �?      A@      @              @      A@              <@      6@      <@      1@              @      <@      &@      "@       @      "@                       @      3@      "@              @      3@      @      @       @               @      @              .@      @      .@                      @              @      1@      ;@      @      7@      @      *@      @      @      @              @      @      @       @       @      �?              �?       @              �?      �?              �?      �?              �?      @      �?      �?              �?      �?                      @              @              $@      $@      @      @              @      @      @               @      @       @      �?       @                      �?              @     �p@      0@     �p@      &@     �j@      �?     �h@              3@      �?      @      �?              �?      @              *@             �H@      $@      4@       @      4@      �?      3@              �?      �?              �?      �?                      �?      =@       @      =@      @      1@              (@      @      (@      @      @      @      @      @      @              �?      @              @      �?               @              @                       @               @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK텔h~�B�3         �       
             �?>���i��?2           ��@       I                   �a@
�e4���?C            �@       6       	          pff�?Dcq1��?�            0x@       5                    �R@$�� ���?�            �m@       0                    �?p�)_�5�?�            �m@              	          ����?Ld����?`            �c@       
                    �?�O4R���?#            �J@       	                   Pf@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        !             I@                           �?t�n_Y��?=             Z@                           �G@�n_Y�K�?
             *@������������������������       �                      @                          �W@���!pc�?	             &@������������������������       �                     @              	          ����?      �?              @                           �?r�q��?             @                          �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @       %                   P`@�θ�?3            �V@                          �a@b�2�tk�?             B@������������������������       �                      @              	          ����?      �?             <@������������������������       �                     @                          Pj@� �	��?             9@������������������������       �                     @                            �?�<ݚ�?             2@������������������������       �                      @!       "                    �?      �?             0@������������������������       �                     $@#       $                   �`@�q�q�?             @������������������������       �                     @������������������������       �                      @&       '                     F@X�;�^o�?            �K@������������������������       �                      @(       )                    `@0��_��?            �J@������������������������       �                     F@*       +                   �`@X�<ݚ�?             "@������������������������       �                     @,       -                    �?�q�q�?             @������������������������       �                     @.       /                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @1       4                   �X@�Fǌ��?1            �S@2       3                    �?��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@������������������������       �        )             P@������������������������       �                      @7       8                   �U@hڛ�ʚ�?]            �b@������������������������       �                     �?9       >                    �?�?�|�?\            �b@:       =                    �?�r����?	             .@;       <                    �O@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     &@?       F                    �R@���%yU�?S            �`@@       E                    �J@�7�	|��?P             `@A       B                   �o@г�wY;�?             A@������������������������       �                     3@C       D                    @J@��S�ۿ?
             .@������������������������       �        	             ,@������������������������       �                     �?������������������������       �        :            �W@G       H                   �p@      �?             @������������������������       �                     @������������������������       �                     �?J       O                   e@�K��&�?T             `@K       L                    �?�nkK�?             7@������������������������       �                     5@M       N       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?P       }                    �?      �?D            �Z@Q       l                    @L@,�|%�v�?6            @U@R       W                    �?ҐϿ<��?$            �N@S       T                   q@�}�+r��?
             3@������������������������       �                     0@U       V                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @X       k                   �a@�G��l��?             E@Y       \                    �?�Gi����?            �B@Z       [                   �e@���!pc�?             &@������������������������       �                      @������������������������       �                     @]       ^                   �m@R�}e�.�?             :@������������������������       �                     *@_       j                    �?��
ц��?             *@`       i                    �?���Q��?             $@a       b                    �?      �?              @������������������������       �                     @c       d                    ]@���Q��?             @������������������������       �                     �?e       h                    �?      �?             @f       g                   �o@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @m       n       
             �?�q�q�?             8@������������������������       �                     �?o       |                    @8����?             7@p       {                    �?���!pc�?             6@q       z                    �?�q�q�?             2@r       w                    �?z�G�z�?
             .@s       t                   �q@�q�q�?             @������������������������       �                     @u       v                    b@�q�q�?             @������������������������       �                      @������������������������       �                     �?x       y                     O@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?~       �                   �d@���N8�?             5@       �                    �?�����H�?             2@������������������������       �                     &@�       �                   �n@����X�?             @�       �                   0d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       	          ����?Ɩ�/���?�             y@�       �                    ]@؇���X�?�             t@�       �                    �?��N`.�?#            �K@�       �                   g@�LQ�1	�?             7@������������������������       �                     "@�       �                   �b@և���X�?             ,@������������������������       �                     @�       �                   �[@؇���X�?             @�       �       	          ����?      �?             @�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?     ��?             @@�       �                    �G@�����H�?             ;@�       �                    �?�z�G��?             $@������������������������       �                     @�       �                    @���Q��?             @�       �                   @[@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     1@������������������������       �                     @�       �                    �?��c+��?�            �p@�       �                    �?�|����?�            `m@�       �                   �X@�Wv���?{             k@�       �                   �V@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �b@0z�(>��?y            �j@�       �                    @L@�X-:oȤ?n             h@������������������������       �        \            �d@�       �                   �h@8�Z$���?             :@������������������������       �                      @�       �                    b@�<ݚ�?             2@�       �       	            �?@�0�!��?
             1@�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                   @`@      �?              @������������������������       �                     @�       �                   @t@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   p`@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                     R@      �?             4@�       �                   �c@r�q��?
             2@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     *@������������������������       �                      @�       �                   �h@�\��N��?             3@������������������������       �                     @�       �                    �?���Q��?             .@�       �                   �p@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   `R@     ��?             @@������������������������       �                     @�       �                   �o@\-��p�?             =@������������������������       �        
             0@�       �       	          @33�?�	j*D�?             *@�       �                    �?���|���?             &@�       �                    �?և���X�?             @�       �                   �r@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?R�����?3             T@�       �                    �?�q����?#            �J@������������������������       �        
             0@�       �       	          ����?��J�fj�?            �B@������������������������       �                     @�       �                   �p@�4�����?             ?@�       �       	          033@��}*_��?             ;@�       �                   �n@��+7��?             7@�       �                    �?��s����?             5@�       �                    �I@�q�q�?             (@������������������������       �                      @�       �                   �_@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     "@������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �Z@�<ݚ�?             ;@������������������������       �        
             2@�       �                    �M@�q�q�?             "@������������������������       �                     @�       �                    �?      �?             @�       �                   Xw@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@      W@     �z@      C@     �u@     �@@     �i@      ?@     �i@      >@     �_@      �?      J@      �?       @      �?                       @              I@      =@     �R@       @      @               @       @      @      @              @      @      @      �?       @      �?       @                      �?      @                       @      5@     �Q@      ,@      6@               @      ,@      ,@      @              &@      ,@      @              @      ,@       @               @      ,@              $@       @      @              @       @              @      H@       @              @      H@              F@      @      @      @               @      @              @       @      �?              �?       @              �?     �S@      �?      ,@      �?                      ,@              P@       @              @      b@      �?              @      b@       @      *@       @       @               @       @                      &@       @     ``@      �?      `@      �?     �@@              3@      �?      ,@              ,@      �?                     �W@      �?      @              @      �?              K@     �R@      �?      6@              5@      �?      �?              �?      �?             �J@     �J@      H@     �B@      D@      5@      2@      �?      0@               @      �?              �?       @              6@      4@      6@      .@      @       @               @      @              3@      @      *@              @      @      @      @      @       @      @              @       @      �?               @       @      �?       @      �?                       @      �?                       @              @              @       @      0@      �?              @      0@      @      0@      @      (@      @      (@       @      @              @       @      �?       @                      �?      �?       @               @      �?              @                      @      �?              @      0@       @      0@              &@       @      @       @      �?       @                      �?              @      @             �s@     �T@     @q@      G@     �B@      2@       @      .@              "@       @      @      @              �?      @      �?      @      �?      �?              �?      �?                       @              @      =@      @      8@      @      @      @      @               @      @      �?      @              @      �?              �?              1@              @             �m@      <@     �j@      5@     �i@      &@      �?       @      �?                       @     �i@      "@     �g@      @     �d@              6@      @       @              ,@      @      ,@      @      $@      �?      @              @      �?      @              �?      �?      �?                      �?      @       @               @      @                      �?      .@      @      .@      @       @      @       @                      @      *@                       @      "@      $@              @      "@      @      @      @      @                      @      @              9@      @              @      9@      @      0@              "@      @      @      @      @      @      @      �?      @                      �?              @      @               @             �E@     �B@     �B@      0@      0@              5@      0@              @      5@      $@      1@      $@      1@      @      1@      @       @      @               @       @       @               @       @              "@                       @              @      @              @      5@              2@      @      @      @              �?      @      �?      �?              �?      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�lBLhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKم�h~�Bx/         x       
             �?��e�B��??           ��@       	                   �a@��k��?I           X�@                          �a@P����?O            �]@������������������������       �        D            @Y@                           �?�t����?             1@������������������������       �        	             ,@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?
       '                    �?���iz�?�            Py@                          �\@�\����?-            �P@������������������������       �                     &@       &       	             @���|���?'            �K@       %                    �?����X�?"            �H@                           �a@�5��
J�?              G@                           �K@�?�'�@�?             C@                            I@�nkK�?             7@������������������������       �        
             .@                           �?      �?              @������������������������       �                     �?                          @_@؇���X�?             @������������������������       �                     @                          Hp@      �?             @������������������������       �                     @������������������������       �                     �?              	          @33�?������?             .@������������������������       �                     @                           �?�8��8��?	             (@������������������������       �                     $@              	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?!       $       	          033�?      �?              @"       #                   �`@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @(       ]                   P`@4�^o�]�?�            0u@)       P                   �b@~���)r�?g            �d@*       +       
             �?f>�cQ�?O            �^@������������������������       �                     *@,       K                    �?6�����?H            @[@-       @                    �?��T|n�?;            �U@.       3                   �Z@���}<S�?/            @Q@/       0                   `_@      �?              @������������������������       �                     @1       2                   `W@      �?             @������������������������       �                     �?������������������������       �                     @4       ?                   �k@�.ߴ#�?)            �N@5       6                   @_@H%u��?             9@������������������������       �                     $@7       >                   �k@z�G�z�?             .@8       9                   �h@؇���X�?
             ,@������������������������       �                     @:       =                    �L@      �?              @;       <                   �j@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     B@A       F                   �a@��.k���?             1@B       E                     N@      �?              @C       D                     K@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @G       J                    ]@�����H�?             "@H       I                   `b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @L       M                    @P@�LQ�1	�?             7@������������������������       �                     3@N       O                    �P@      �?             @������������������������       �                     @������������������������       �                     �?Q       T                    ]@��Hg���?            �F@R       S                   �q@�q�q�?             @������������������������       �                     @������������������������       �                      @U       V       
             �?:�&���?            �C@������������������������       �                     ,@W       X                   0o@ �o_��?             9@������������������������       �                     1@Y       Z                     O@      �?              @������������������������       �                     @[       \       	          833�?      �?              @������������������������       �                     �?������������������������       �                     �?^       a                     E@�Ts�k��?f            �e@_       `                   �i@�q�q�?             @������������������������       �                      @������������������������       �                     �?b       q                    @ps��pй?c             e@c       p                    �?���j�?[            @c@d       e                    a@X�?٥�?<            �Y@������������������������       �        +            @T@f       g                   Pa@�GN�z�?             6@������������������������       �                      @h       i                     L@R���Q�?             4@������������������������       �                     $@j       o                    �?�z�G��?             $@k       l                   �b@���Q��?             @������������������������       �                      @m       n       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                    �I@r       w                   �o@������?             .@s       v                    �?և���X�?             @t       u                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @y       �                    �L@4�ƙ���?�            �x@z       �                    �?TO|?=��?�            �r@{       �       	             @�Aʑ���?�            �p@|       �                   �e@<ASĹ�?�            �p@}       ~                    �?�q�q�?             >@������������������������       �                     @       �                    �?r�q��?             8@�       �                   �X@���N8�?             5@������������������������       �                     �?������������������������       �                     4@������������������������       �                     @�       �                    �?86��Z�?�            �m@�       �                   �b@d}h���?"             L@�       �                   �b@8�Z$���?!             J@������������������������       �                     1@�       �                     B@4�2%ޑ�?            �A@������������������������       �                     �?�       �                    �E@H�V�e��?             A@������������������������       �                     &@�       �                   �f@8����?             7@�       �                    @J@��S���?             .@�       �                    �?�z�G��?             $@������������������������       �                      @�       �                    b@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    @L@�rǬ鰠?q            �f@�       �                   @n@�E�����?p            �f@������������������������       �        ?            �X@�       �                     G@��Y��]�?1            �T@������������������������       �                    �F@�       �                   pn@@-�_ .�?            �B@������������������������       �                     �?�       �                    �?������?             B@�       �                   0q@؇���X�?             @������������������������       �                     @�       �                    @J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     =@������������������������       �                     �?������������������������       �                     @�       �                    �?��}*_��?             ;@�       �                   @[@�θ�?	             *@������������������������       �                     "@�       �                    �H@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             ,@�       �       	          ����?D�]�+��?=            �X@�       �                   @\@�j�'�=�?*            �P@�       �                   �Z@���|���?             &@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �b@�rF���?"            �K@�       �                   `_@(;L]n�?             >@�       �                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     4@�       �       	          pff�?� �	��?             9@�       �                    �?�G��l��?             5@�       �                    _@�<ݚ�?             "@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                     O@�q�q�?             (@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                    s@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                     P@      �?             @@�       �                    @N@8�Z$���?             :@�       �                    �?�q�q�?             (@������������������������       �                     @�       �                   �a@      �?              @�       �                    �?�q�q�?             @�       �       	          033�?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     ,@�       �                   �b@�q�q�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�b�     h�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@      Y@     pz@       @      ]@             @Y@       @      .@              ,@       @      �?       @                      �?     �X@     0s@     �A@      ?@              &@     �A@      4@     �A@      ,@     �A@      &@     �@@      @      6@      �?      .@              @      �?      �?              @      �?      @              @      �?      @                      �?      &@      @              @      &@      �?      $@              �?      �?      �?                      �?       @      @      �?      @      �?                      @      �?                      @              @     �O@     @q@      J@     �\@      2@      Z@              *@      2@     �V@      .@     �Q@      @     �O@      @      @              @      @      �?              �?      @              @      M@      @      6@              $@      @      (@       @      (@              @       @      @       @      @       @                      @               @      �?                      B@      "@       @      �?      @      �?      @              @      �?                      @       @      �?      @      �?      @                      �?      @              @      4@              3@      @      �?      @                      �?      A@      &@       @      @              @       @              @@      @      ,@              2@      @      1@              �?      @              @      �?      �?              �?      �?              &@      d@       @      �?       @                      �?      "@      d@      @     �b@      @     �X@             @T@      @      1@       @              @      1@              $@      @      @      @       @       @              �?       @      �?                       @              @             �I@      @      &@      @      @      @      �?      @                      �?               @               @     �s@     @T@     0p@      C@     @n@      <@     @n@      9@      4@      $@              @      4@      @      4@      �?              �?      4@                      @     �k@      .@      F@      (@      F@       @      1@              ;@       @              �?      ;@      @      &@              0@      @       @      @      @      @       @              �?      @              @      �?              @               @                      @     @f@      @     @f@       @     �X@              T@       @     �F@             �A@       @              �?     �A@      �?      @      �?      @              �?      �?      �?                      �?      =@                      �?              @      1@      $@      @      $@              "@      @      �?              �?      @              ,@             �K@     �E@     �G@      3@      @      @              @      @       @      @                       @     �E@      (@      =@      �?      "@      �?              �?      "@              4@              ,@      &@      $@      &@       @      @       @      @       @                      @              @       @      @      @      �?              �?      @              �?      @      �?                      @      @               @      8@      @      6@      @       @              @      @      @       @      @       @       @               @       @                       @       @                      ,@      @       @      �?       @      �?                       @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��V-hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK߅�h~�B�0         �                    �?>���i��?L           ��@       K                    �?�ԍ�LN�?>           �~@       @                    �?��k��&�?�             j@       =       	          ����?Vǃ���?Y            �a@       6                    �?     ��?O             `@       	                   @E@o�����?F             ]@                          pb@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @
       )                   �_@������?>            �Y@       &                   Xr@���b���?!            �L@                          d@ҳ�wY;�?            �I@              
             �?��Q���?             D@                          �p@����X�?             ,@                           _@�C��2(�?             &@������������������������       �                     @                          �d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                          �a@R�}e�.�?             :@                           `P@؇���X�?             @������������������������       �                     @������������������������       �                     �?                           �?�}�+r��?             3@������������������������       �                     �?������������������������       �                     2@                          `i@���|���?             &@������������������������       �                      @       %                    _@�<ݚ�?             "@                           `]@      �?              @������������������������       �                     @!       "                    �?      �?             @������������������������       �                     �?#       $                    �B@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?'       (                   ``@r�q��?             @������������������������       �                     �?������������������������       �                     @*       1       
             �?��+7��?             G@+       ,       	          ����?������?
             .@������������������������       �                     @-       .                    �?X�<ݚ�?             "@������������������������       �                     @/       0                   �_@z�G�z�?             @������������������������       �                     �?������������������������       �                     @2       5                    �D@�g�y��?             ?@3       4                   @b@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     8@7       8                    @K@�8��8��?	             (@������������������������       �                     @9       <                   �^@؇���X�?             @:       ;                    @L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @>       ?       
             �?$�q-�?
             *@������������������������       �        	             (@������������������������       �                     �?A       B                   Pj@t�U����?)            �P@������������������������       �                    �H@C       D                   n@X�<ݚ�?             2@������������������������       �                     @E       F                   @Y@�q�q�?	             .@������������������������       �                     @G       H                    �?�C��2(�?             &@������������������������       �                     @I       J                   u@      �?              @������������������������       �                     @������������������������       �                     �?L       o       	          ����?x�}b~|�?�            �q@M       b                    �?�4�M�f�?D            �Y@N       S                    a@R���Q�?5             T@O       P                   �s@      �?             @@������������������������       �                     >@Q       R                    �?      �?              @������������������������       �                     �?������������������������       �                     �?T       U                   �j@�q�q��?             H@������������������������       �        
             0@V       ]                    @I@     ��?             @@W       X                   �\@r�q��?             (@������������������������       �                     �?Y       Z                    @H@�C��2(�?             &@������������������������       �                     "@[       \       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?^       a                     L@P���Q�?             4@_       `                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     1@c       n                   �e@�X����?             6@d       m                    �N@      �?             4@e       f                   `X@�q�q�?	             (@������������������������       �                      @g       l                    @N@�z�G��?             $@h       i                   �]@�<ݚ�?             "@������������������������       �                     �?j       k       
             �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @p       u                    �?�]0��<�?x            �f@q       r                   @a@R���Q�?             4@������������������������       �                     $@s       t                   Pi@�z�G��?             $@������������������������       �                     @������������������������       �                     @v       w                   �U@�\����?l            `d@������������������������       �                     �?x       }       
             �? �)���?k            @d@y       z       	          033@ ���?^             b@������������������������       �        I            @\@{       |                   �Z@      �?             @@������������������������       �                     �?������������������������       �                     ?@~                           c@�IєX�?             1@������������������������       �                     0@������������������������       �                     �?�       �                   `@��A��?           �z@�       �       
             �?$ޗQ��?@            �Y@�       �                    �?��v����?(            �P@�       �                    �?�û��|�?             7@�       �                     P@      �?              @�       �       	          ����?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?z�G�z�?	             .@�       �                   `X@�z�G��?             $@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    `Q@؇���X�?             @������������������������       �                     @�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     F@�       �                     P@�#-���?            �A@�       �                    Y@      �?             @@������������������������       �                     �?������������������������       �                     ?@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       
             �?@�0�!��?�            0t@�       �                    �?��
P��??            @Z@�       �                   �_@�q�q�?            �@@������������������������       �                     (@�       �                    �?�G��l��?             5@�       �       	          ����?j���� �?
             1@�       �                    �H@�q�q�?             "@������������������������       �                      @�       �                   �a@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                   �g@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       	          pff�?P��E��?,             R@�       �                    f@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                   �o@N1���?&            �N@�       �                   b@D�n�3�?             C@�       �                   0m@؇���X�?             ,@�       �                   pa@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?�       �                   �m@�q�q�?             8@�       �                   �a@�d�����?             3@�       �                   �c@     ��?             0@������������������������       �                     "@�       �                   @d@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �b@�q�q�?             @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       
             �?��+7��?             7@������������������������       �                     @�       �                    �?R���Q�?             4@�       �                    @H@�q�q�?             "@������������������������       �                     @�       �                    �?      �?             @�       �                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�       �                    @`���˛?�            @k@�       �                    �?`�LVXz�?�            �h@�       �                    �O@����7�?r             f@�       �                   @g@�����?o            �e@������������������������       �        n            �e@������������������������       �                     �?�       �                   Pc@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     5@�       �                   �j@P���Q�?             4@�       �                   �`@�����H�?             "@�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@      Z@     Px@     �S@      `@     �Q@     �Q@     �Q@      M@     �M@     �L@       @      &@              &@       @             �L@      G@      7@      A@      2@     �@@      &@      =@      @      $@      �?      $@              @      �?      @      �?                      @      @              @      3@      @      �?      @                      �?      �?      2@      �?                      2@      @      @               @      @       @      @      �?      @              @      �?      �?               @      �?       @                      �?              �?      @      �?              �?      @              A@      (@      @      &@              @      @      @              @      @      �?              �?      @              >@      �?      @      �?      @                      �?      8@              &@      �?      @              @      �?       @      �?              �?       @              @              �?      (@              (@      �?               @     �M@             �H@       @      $@      @              @      $@      @              �?      $@              @      �?      @              @      �?              9@     @p@      3@     �T@      (@      Q@      �?      ?@              >@      �?      �?      �?                      �?      &@     �B@              0@      &@      5@      $@       @              �?      $@      �?      "@              �?      �?              �?      �?              �?      3@      �?       @      �?                       @              1@      @      .@      @      .@      @      @       @              @      @       @      @      �?              �?      @              @      �?              �?                       @       @              @      f@      @      1@              $@      @      @      @                      @      @      d@      �?               @      d@      �?      b@             @\@      �?      ?@      �?                      ?@      �?      0@              0@      �?             0s@     �]@     �D@     �N@      "@      M@      "@      ,@      @       @       @       @       @                       @      @              @      (@      @      @       @      �?       @                      �?      �?      @              @      �?       @               @      �?                      @              F@      @@      @      ?@      �?              �?      ?@              �?       @      �?                       @     �p@     �L@     �I@      K@      6@      &@      (@              $@      &@      $@      @      @      @       @              �?      @              @      �?              @      �?              �?      @                      @      =@     �E@      �?      $@              $@      �?              <@     �@@      6@      0@      (@       @      (@      �?              �?      (@                      �?      $@      ,@      @      ,@      @      *@              "@      @      @      @                      @       @      �?      �?              �?      �?              �?      �?              @              @      1@      @              @      1@      @      @              @      @      �?       @      �?       @                      �?      �?                      &@     �j@      @     �h@       @     �e@       @     �e@      �?     �e@                      �?      @      �?      @                      �?      5@              3@      �?       @      �?       @      �?       @                      �?      @              &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��@hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM'hwh(h+K ��h-��R�(KM'��h~�B�@         �                    �?��t�?>           ��@       1                    �?�Q�N��?T           ��@       (                    �?��-*�?b            @b@                           �?��ϻ�r�?X            ``@                           �?�!���?             A@                           b@j���� �?             1@������������������������       �                      @       	                   pc@�q�q�?
             .@������������������������       �                     @
                           `@      �?             $@������������������������       �                     @              	          `ff�?����X�?             @                          �p@���Q��?             @������������������������       �                     �?              
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @              
             �?�IєX�?
             1@                          �R@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@                          `X@h�a��?B            @X@������������������������       �                     �?       %       
             �? �q�q�?A             X@                          �b@ �Cc}�?             <@������������������������       �                     &@       "                   hq@@�0�!��?             1@                            L@$�q-�?             *@������������������������       �                     $@        !                    �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @#       $                   �q@      �?             @������������������������       �                      @������������������������       �                      @&       '                     R@ ��ʻ��?/             Q@������������������������       �        .            �P@������������������������       �                     �?)       ,                    �?���Q��?
             .@*       +                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @-       0       	          ����?z�G�z�?             $@.       /       
             �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     �?2       Y                   @E@�a����?�            �x@3       J       
             �?"�W1��?2            �T@4       ;       	          ����?���c���?!             J@5       :                   �X@`2U0*��?             9@6       9                    �?      �?             @7       8                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     5@<       A                    �?�<ݚ�?             ;@=       @       
             �?�����H�?
             2@>       ?                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     (@B       C                   �_@X�<ݚ�?             "@������������������������       �                      @D       E                    �I@և���X�?             @������������������������       �                     �?F       G                    �P@�q�q�?             @������������������������       �                     @H       I       	          hff @�q�q�?             @������������������������       �                     �?������������������������       �                      @K       V                     P@�q�q�?             >@L       Q                   �`@��<b���?             7@M       N                   �W@և���X�?             @������������������������       �                      @O       P       	          ����?z�G�z�?             @������������������������       �                     @������������������������       �                     �?R       S                    �?      �?             0@������������������������       �                     &@T       U                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?W       X       	          `ff�?����X�?             @������������������������       �                     @������������������������       �                      @Z       �       	          ����?n�����?�            �s@[       h                   @]@    ���?�             p@\       g                   @f@r�q��?             H@]       ^                    �?�&!��?            �E@������������������������       �                     @_       `       
             �?)O���?             B@������������������������       �                     0@a       b                    @G@R���Q�?             4@������������������������       �                      @c       f                    �G@      �?             (@d       e                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @i       �       	          833�?��ջ�A�?�             j@j       �                   �f@�S����?`             c@k       �                    @T;���?Y            �a@l       �                    �?��v����?U            �`@m       x                   �a@�^����?J            �]@n       w                    �O@`�H�/��?>            �Y@o       v                   a@��T�u��?=            @Y@p       s                   �`@��v����?*            �P@q       r       
             �?Xny��?%            �N@������������������������       �                     @������������������������       �                      K@t       u                   0q@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     A@������������������������       �                     �?y       �                     M@      �?             0@z                          `z@؇���X�?
             ,@{       ~                    �D@$�q-�?	             *@|       }                   �b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             0@�       �                    �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?���Q��?             @�       �                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                     O@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                   pa@Dc}h��?              L@�       �                   Pd@ףp=
�?             4@������������������������       �        	             2@������������������������       �                      @�       �       
             �?�q�q�?             B@�       �                    �?�G�z��?             4@�       �                   @c@�����H�?             "@�       �                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          833�?���!pc�?             &@������������������������       �                      @�       �                    �?�����H�?             "@�       �                    `P@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             0@������������������������       �                      @�       �       	          pff�?؇���X�?             ,@�       �                    a@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@�       �       
             �?$gv&��?$            �M@�       �       
             �?ףp=
�?             I@�       �                     O@և���X�?             @������������������������       �                     @������������������������       �                     @�       �       	          `ff�? �#�Ѵ�?            �E@�       �       	          `ff�?�����H�?             "@������������������������       �                     @�       �                   p@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �n@г�wY;�?             A@������������������������       �                     9@�       �                    �?�����H�?             "@������������������������       �                     @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   (p@�<ݚ�?             "@������������������������       �                     @�       �                    �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @�                         �b@�J�4�?�            pw@�       �       
             �?���H��?�             u@�       �                   �]@l������?�            �r@�       �                    �?��Y��]�?O            �^@�       �                    �?�E�����?:            �V@�       �       	          433�? ��ʻ��?/             Q@�       �                   �Y@�IєX�?             1@������������������������       �                     &@�       �       	          ����?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        $            �I@������������������������       �                     6@�       �                    �?�FVQ&�?            �@@�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?h�����?             <@�       �                   `c@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     6@�       �                   �Z@H%u��?k            �e@�       �                   `l@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�       �                   �s@�5U��K�?g            �d@�       �                   �b@�.(�i��?_            �b@�       �                    �?(;L]n�?K             ^@�       �                   �`@"pc�
�?             &@�       �                    �N@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       	          033�?����q�?F            @[@������������������������       �        "            �J@�       �       	          `ff�?h�����?$             L@�       �                    @�<ݚ�?             "@�       �                   �i@      �?              @�       �                     G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                    �G@�       �                   �a@�n`���?             ?@�       �                    �N@���!pc�?             6@�       �       	             �?      �?             0@�       �                     M@      �?             (@�       �       	             �?      �?              @������������������������       �                      @�       �                     I@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                   ht@���Q��?             .@������������������������       �                     @�       �                   �u@ףp=
�?             $@������������������������       �                     @�       �                    @L@      �?             @������������������������       �                     @������������������������       �                     �?                          �N@D�n�3�?             C@            	             �?|��?���?             ;@                         �?ףp=
�?             $@                         @I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                         �?�t����?             1@                        �^@z�G�z�?             .@	      
      	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                         c@�8��8��?
             (@������������������������       �                     $@                         `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                        �l@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @            
             �?Hث3���?            �C@            	          ����?�E��ӭ�?
             2@������������������������       �                     @                         c@@4և���?             ,@                         �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@      &                   �?����X�?             5@                         �J@���Q��?             $@������������������������       �                     @       !                   _@�q�q�?             @������������������������       �                     �?"      #                   a@z�G�z�?             @������������������������       �                      @$      %                   d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KM'KK��h_�Bp       �x@     8�@     0u@     �i@     @^@      9@     �\@      0@      7@      &@      @      $@       @              @      $@              @      @      @      @               @      @       @      @      �?              �?      @      �?                      @               @      0@      �?      @      �?              �?      @              *@              W@      @              �?      W@      @      9@      @      &@              ,@      @      (@      �?      $@               @      �?              �?       @               @       @               @       @             �P@      �?     �P@                      �?      @      "@      @      �?              �?      @               @       @       @      @              @       @                      �?     @k@     `f@      1@     @P@      @     �F@      �?      8@      �?      @      �?       @               @      �?                      �?              5@      @      5@       @      0@       @      @              @       @                      (@      @      @               @      @      @              �?      @       @      @              �?       @      �?                       @      $@      4@      @      2@      @      @               @      @      �?      @                      �?      �?      .@              &@      �?      @              @      �?              @       @      @                       @      i@     �\@     �g@     �P@      6@      :@      1@      :@              @      1@      3@              0@      1@      @       @              "@      @      �?      @      �?                      @       @              @             �d@     �D@      `@      8@     �]@      8@      ]@      2@      Z@      ,@      W@      $@      W@      "@      M@      "@      K@      @              @      K@              @       @      @                       @      A@                      �?      (@      @      (@       @      (@      �?      @      �?      @                      �?      "@                      �?               @      (@      @      $@      �?      $@                      �?       @      @       @      �?       @                      �?               @      @      @              @      @              "@             �C@      1@      2@       @      2@                       @      5@      .@      "@      &@      �?       @      �?       @               @      �?                      @       @      @               @       @      �?      @      �?      @                      �?       @              (@      @               @      (@       @      @       @               @      @              "@              (@     �G@      @     �F@      @      @              @      @               @     �D@      �?       @              @      �?      �?      �?                      �?      �?     �@@              9@      �?       @              @      �?      �?      �?                      �?      @       @      @              �?       @      �?                       @      N@     �s@      D@     �r@      8@      q@      @      ^@      �?     @V@      �?     �P@      �?      0@              &@      �?      @              @      �?                     �I@              6@       @      ?@      �?      @              @      �?              �?      ;@      �?      @              @      �?                      6@      5@     @c@      @      @      @                      @      0@     �b@      $@     �a@      @      ]@       @      "@       @      @       @                      @              @       @     �Z@             �J@       @      K@       @      @      �?      @      �?      �?              �?      �?                      @      �?                     �G@      @      9@      @      0@      @      $@      @      @       @      @               @       @      @       @                      @      @                      @              @              "@      @      "@      @              �?      "@              @      �?      @              @      �?              0@      6@      ,@      *@      "@      �?       @      �?              �?       @              @              @      (@      @      (@       @      �?              �?       @              �?      &@              $@      �?      �?      �?                      �?       @               @      "@              "@       @              4@      3@      @      *@      @              �?      *@      �?      @      �?                      @              $@      .@      @      @      @              @      @       @              �?      @      �?       @               @      �?              �?       @              &@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJۋ�<hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B(5         �       
             �?:���sQ�?;           ��@       M                    �?p��#�?B           @@       (                   �b@@ �h�\�?�            @i@              	          ����?<���D�?W            �`@                          �X@���#�İ?%            �M@                          `Z@�C��2(�?             &@       
                    �?      �?              @       	                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           �E@@��8��?             H@                           �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     E@              	          pff�?��W��?2            @R@                          �a@r�q��?             8@                           b@d}h���?             ,@������������������������       �                     $@                          �b@      �?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     $@       %                    �Q@��<D�m�?             �H@                            �?�nkK�?             G@                          @_@r�q��?             @������������������������       �                     �?������������������������       �                     @!       "                   �b@�(\����?             D@������������������������       �                    �B@#       $                   Pd@�q�q�?             @������������������������       �                     �?������������������������       �                      @&       '                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @)       0                    �?B� ��?.            �Q@*       /                    b@�<ݚ�?             ;@+       ,                   �Q@      �?             8@������������������������       �                     �?-       .       	          ���@���}<S�?             7@������������������������       �                     5@������������������������       �                      @������������������������       �                     @1       6                    �D@�K��&�?            �E@2       3                    �?      �?              @������������������������       �                     @4       5                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @7       B                    �?��
P��?            �A@8       A                   �`@p�ݯ��?             3@9       >                   8p@z�G�z�?	             .@:       ;                   �j@�C��2(�?             &@������������������������       �                     @<       =                   �]@r�q��?             @������������������������       �                     �?������������������������       �                     @?       @                   Pr@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @C       F                   0m@     ��?             0@D       E       	             @�����H�?             "@������������������������       �                      @������������������������       �                     �?G       H                   `]@և���X�?             @������������������������       �                     �?I       L                   pb@�q�q�?             @J       K                   �c@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?N       O                   Pe@Ъ�U��?�            �r@������������������������       �        -            @Q@P       U                   �f@��Q�Vz�?�            �l@Q       R                   �a@և���X�?             @������������������������       �                     @S       T                   �e@      �?             @������������������������       �                     �?������������������������       �                     @V       }                    �?,N�_� �?�            �k@W       X                   �Z@�f�?g            `d@������������������������       �                      @Y       z                    �R@@�#����?e             d@Z       w                    @0G���ջ?c            �c@[       p                   �m@�kb97�?a            @c@\       e                   @^@ ����?&            @P@]       ^                    Y@     ��?
             0@������������������������       �                     �?_       b                   0i@�r����?	             .@`       a                   ph@      �?              @������������������������       �                     �?������������������������       �                     �?c       d                   �b@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?f       i                    @H@Hm_!'1�?            �H@g       h                   �k@      �?             @������������������������       �                     �?������������������������       �                     @j       o                   �[@����?�?            �F@k       n       	             �?�����H�?             "@l       m       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     B@q       v                   0q@ }�Я��?;            @V@r       s       	          `ff�? ���J��?            �C@������������������������       �                     8@t       u                   `b@��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �        "             I@x       y                    @Q@      �?              @������������������������       �                     �?������������������������       �                     �?{       |       	             @���Q��?             @������������������������       �                     @������������������������       �                      @~       �                   �_@P����?$            �M@       �                    �?z�G�z�?             @�       �                   �^@      �?             @�       �                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     K@�       �                    �?b��K�?�             z@�       �                   @E@������?�            `v@�       �       	          `ff�?�KM�]�?             C@�       �                   �X@���y4F�?             3@������������������������       �                     @�       �                    �?�	j*D�?
             *@�       �                    �N@z�G�z�?             $@�       �                   `\@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             3@�       �                    �?(\����?�             t@�       �                    @N@�����?5            �U@�       �                    @J@R���Q�?0             T@�       �                   �a@���c�H�?!            �H@������������������������       �                     ,@�       �                    �I@">�֕�?            �A@�       �                    �?�������?             >@�       �                   0j@�eP*L��?             &@������������������������       �                     @�       �                   pm@      �?              @������������������������       �                     @�       �                   �c@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   pf@�}�+r��?             3@������������������������       �        	             0@�       �                   �f@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   @Z@�g�y��?             ?@�       �                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     <@�       �       	          `ff�?����X�?             @�       �                   �b@r�q��?             @�       �                   @n@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �g@�!��?�             m@�       �                    �?��[B��?�             m@�       �                    @L@��� ��?             ?@������������������������       �        	             .@�       �                    �?      �?
             0@�       �                   pb@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   `_@8�Z$���?             *@�       �                   `Z@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@�       �                    @L@�/��5�?z             i@�       �                    �G@�Sa��?c            �d@�       �                    �?x�G�z�?0             T@������������������������       �                     >@�       �                    @G@ "��u�?             I@������������������������       �                     G@�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        3            �U@�       �                    �L@�t����?             A@�       �                    �?���Q��?             @�       �       	          @33�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                     P@ 	��p�?             =@�       �                    �O@�t����?             1@�       �                    @��S�ۿ?
             .@������������������������       �        	             ,@������������������������       �                     �?�       �                   @t@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?�       �                   `d@�0u��A�?              N@�       �                    �?�-���?             I@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    @L@"pc�
�?             F@�       �                    @I@     ��?	             0@������������������������       �                      @�       �                    @J@      �?              @�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	          ����?h�����?             <@�       �                    �N@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     7@������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B0       �x@     p�@     �R@     �z@     �K@     `b@      0@      ]@       @     �L@      �?      $@      �?      @      �?      @              @      �?                      @              @      �?     �G@      �?      @              @      �?                      E@      ,@     �M@      &@      *@      &@      @      $@              �?      @      �?      �?              �?      �?                       @              $@      @      G@       @      F@      �?      @      �?                      @      �?     �C@             �B@      �?       @      �?                       @      �?       @      �?                       @     �C@      ?@      5@      @      5@      @              �?      5@       @      5@                       @              @      2@      9@      �?      @              @      �?       @      �?                       @      1@      2@      (@      @      (@      @      $@      �?      @              @      �?              �?      @               @       @               @       @                      @      @      &@      �?       @               @      �?              @      @              �?      @       @      @      �?              �?      @                      �?      3@     pq@             @Q@      3@     @j@      @      @      @              �?      @      �?                      @      .@     �i@      ,@     �b@       @              (@     �b@      "@     `b@       @     @b@      @      M@      @      *@      �?               @      *@      �?      �?              �?      �?              �?      (@              (@      �?              @     �F@      @      �?              �?      @              �?      F@      �?       @      �?       @               @      �?                      @              B@      �?      V@      �?      C@              8@      �?      ,@              ,@      �?                      I@      �?      �?      �?                      �?      @       @      @                       @      �?      M@      �?      @      �?      @      �?      �?              �?      �?                       @              �?              K@     �s@      Y@     pr@     �O@      @      A@      @      .@              @      @      "@       @       @      �?       @      �?                       @      �?               @      �?      �?              �?      �?      �?                      �?              3@     0r@      =@     �Q@      1@      Q@      (@      C@      &@      ,@              8@      &@      7@      @      @      @              @      @      @      @               @      @              @       @              2@      �?      0@               @      �?              �?       @              �?      @              @      �?              >@      �?       @      �?       @                      �?      <@               @      @      �?      @      �?       @      �?                       @              @      �?             �k@      (@     �k@      &@      ;@      @      .@              (@      @      �?       @      �?                       @      &@       @       @       @       @                       @      "@             @h@      @     �d@      @     @S@      @      >@             �G@      @      G@              �?      @              @      �?             �U@              >@      @      @       @      �?       @      �?                       @       @              ;@       @      .@       @      ,@      �?      ,@                      �?      �?      �?      �?                      �?      (@                      �?      7@     �B@      *@     �B@      @      �?      @                      �?       @      B@      @      "@               @      @      �?      @      �?      @                      �?      @              �?      ;@      �?      @      �?                      @              7@      $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��ehG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B�4         �                    �?�	����?E           ��@                           _@���'�?R           8�@              
             �?��A��?9             W@                           �?����˵�?&            �M@������������������������       �                     @                           �? �h�7W�?#            �J@                          �X@�S����?
             3@������������������������       �                     �?	                           �?�����H�?	             2@
                            O@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     &@������������������������       �                     A@                           �N@:ɨ��?            �@@                           \@���B���?             :@              	          `ff�?      �?              @������������������������       �                     @������������������������       �                     @                          @E@�����H�?
             2@������������������������       �        	             0@������������������������       �                      @                           �?����X�?             @������������������������       �                     @������������������������       �                      @       Y       
             �?N\d����?           �|@       N                    �?�lg����?W             `@       C                   @a@�ʻ����?D            �Y@       (       	          ����?��%��?0            �R@       !                    �?@�0�!��?             1@                            �I@      �?              @������������������������       �                     �?������������������������       �                     �?"       '                   �i@�r����?             .@#       $                   `@����X�?             @������������������������       �                     @%       &                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @)       @                   q@���dQ'�?"            �L@*       ;                   @^@ �o_��?             I@+       2                   �a@      �?             8@,       -       	          ����?�	j*D�?             *@������������������������       �                      @.       /                    �?"pc�
�?             &@������������������������       �                     �?0       1                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@3       4                     D@���!pc�?             &@������������������������       �                     �?5       :                    �L@z�G�z�?             $@6       9                   �\@�����H�?             "@7       8                     G@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?<       ?                    �?$�q-�?             :@=       >                     L@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �        
             4@A       B                    �F@؇���X�?             @������������������������       �                     �?������������������������       �                     @D       I                    @�>4և��?             <@E       F                   �x@      �?             8@������������������������       �                     2@G       H                   �a@      �?             @������������������������       �                     @������������������������       �                     @J       K       
             �?      �?             @������������������������       �                     �?L       M                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @O       X                   �x@�����H�?             ;@P       S                   �_@$�q-�?             :@Q       R                    �?      �?              @������������������������       �                     �?������������������������       �                     �?T       U                     Q@ �q�q�?             8@������������������������       �                     4@V       W                   �]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?Z       �                   @g@�FVQ&�?�            �t@[       �       	             @��8=��?�            �t@\       k                    �?hǓ��;�?�            pt@]       j                    �?؇���X�?#             L@^       e                   �q@�ՙ/�?             5@_       b       	          @33�?�θ�?             *@`       a                   g@�����H�?             "@������������������������       �                     �?������������������������       �                      @c       d                   �a@      �?             @������������������������       �                      @������������������������       �                      @f       i                    d@      �?              @g       h                    @I@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                    �A@l       m                   �b@8M��ap�?�            �p@������������������������       �        Q            �`@n       �                    @���.�6�?L            @a@o       x                    �?�5[|/��?H            �`@p       q                    �?��s����?
             5@������������������������       �                     @r       w                   �m@������?             1@s       v                    �G@z�G�z�?             @t       u                   l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@y       z                   c@�?�|�?>            �[@������������������������       �                      @{       �                    �?��wڝ�?=            @[@|       }                    �O@�E�����?3            �V@������������������������       �        0             U@~                           `P@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             3@�       �                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �Z@�	>�p��?�            �v@�       �       	          ����?�eP*L��?             &@������������������������       �                      @�       �                   0a@�q�q�?             "@������������������������       �                     @�       �                   `l@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �b@�+I�9��?�            @v@�       �                    @���)���?�            @t@�       �                    �?\���(�?�             t@�       �                    �J@���y4F�?             C@�       �                    �I@      �?	             ,@�       �                    @I@�z�G��?             $@�       �       	             �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �? �q�q�?             8@������������������������       �        	             1@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?=QcG��?�            �q@�       �                    �R@�0��%�?�            p@�       �                    �N@@�)�n�?�            �o@�       �                    �?�ȉo(��?z            �f@�       �                   �[@�g�y��?i            `c@�       �                    �?�t����?	             1@������������������������       �                     .@������������������������       �                      @�       �                   �[@��<b�ƥ?`            @a@�       �                    @K@l��\��?             A@������������������������       �                     0@�       �                   ph@r�q��?             2@������������������������       �                     "@�       �                   �a@�q�q�?             "@�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        E             Z@�       �       
             �?�����H�?             ;@������������������������       �                     @�       �                   �e@�LQ�1	�?             7@�       �                    �?�C��2(�?             6@�       �                    �L@�r����?	             .@������������������������       �                     $@�       �                   �`@���Q��?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    �? �й���?0            @R@�       �                   (p@�Ń��̧?             E@������������������������       �                    �@@�       �                   �Z@�����H�?             "@�       �       	          ��� @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     ?@�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?`�Q��?             9@�       �                    �?�q�q�?             @������������������������       �                      @�       �                   �Z@      �?             @������������������������       �                     �?�       �                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          ����?���y4F�?             3@������������������������       �                     @�       �                    @L@�	j*D�?	             *@������������������������       �                      @�       �                   `U@"pc�
�?             &@�       �                   �`@���Q��?             @�       �       	          033�?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @L@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?     ��?             @@�       �                    q@r�q��?             8@�       �                    �?�X�<ݺ?             2@�       �       	          433�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             .@�       �                   `q@      �?             @������������������������       �                      @�       �                   �^@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @      �?              @������������������������       �                     @�       �                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?�t�b��"     h�h(h+K ��h-��R�(KK�KK��h_�B        z@     `@     0w@     �f@      *@     �S@      @      L@              @      @      I@      @      0@      �?               @      0@       @      @              @       @                      &@              A@      $@      7@      @      5@      @      @      @                      @       @      0@              0@       @              @       @      @                       @     `v@     @Y@      H@     @T@     �F@     �L@      D@      A@      @      ,@      �?      �?      �?                      �?       @      *@       @      @              @       @      �?              �?       @                       @     �B@      4@      B@      ,@      (@      (@      @      "@       @               @      "@      �?              �?      "@      �?                      "@       @      @              �?       @       @       @      �?       @      �?       @                      �?      @                      �?      8@       @      @       @               @      @              4@              �?      @      �?                      @      @      7@      @      5@              2@      @      @      @                      @       @       @      �?              �?       @      �?                       @      @      8@       @      8@      �?      �?      �?                      �?      �?      7@              4@      �?      @              @      �?              �?             `s@      4@     `s@      2@     `s@      1@      H@       @      *@       @      $@      @       @      �?              �?       @               @       @       @                       @      @      @      @      �?              �?      @                      @     �A@             `p@      "@     �`@              `@      "@     @_@      @      1@      @      @              *@      @      �?      @      �?      �?              �?      �?                      @      (@              [@      @               @      [@      �?     @V@      �?      U@              @      �?              �?      @              3@              @       @               @      @                      �?               @     �F@      t@      @      @       @              @      @              @      @       @      @                       @      D@     �s@      =@     pr@      :@     `r@       @      >@      @      @      @      @      @      @      @                      @              @      @              �?      7@              1@      �?      @              @      �?              2@     �p@      $@     �n@      "@     �n@       @     �e@      @     �b@       @      .@              .@       @              @     �`@      @      ?@              0@      @      .@              "@      @      @      @      �?      @                      �?              @              Z@      @      8@              @      @      4@       @      4@       @      *@              $@       @      @      �?              �?      @              @      �?                      @      �?              �?      R@      �?     �D@             �@@      �?       @      �?      �?      �?                      �?              @              ?@      �?      �?              �?      �?               @      1@      @       @       @               @       @              �?       @      �?       @                      �?      @      .@              @      @      "@       @               @      "@       @      @      �?      @              @      �?              �?                      @      @      �?      @                      �?      &@      5@      @      4@      �?      1@      �?       @      �?                       @              .@      @      @       @              �?      @      �?                      @      @      �?      @              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�;�vhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�7         x       	          ����?�~8�e�?9           ��@       5       
             �?���@�?"           �}@                           �?H�z�'�?]             d@                           �?      �?             @@                           d@������?             ;@                          �q@z�G�z�?             9@                           �?�LQ�1	�?             7@       	                   �Q@�C��2(�?             6@������������������������       �                     �?
                           �?���N8�?
             5@                           �?      �?              @                          Po@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     *@������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @                            �?     ��?K             `@                          �_@*;L]n�?             >@������������������������       �                     &@              	          ����?�����?
             3@                          �l@z�G�z�?             .@                           @K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@                           �?      �?             @������������������������       �                     @������������������������       �                     �?!       $       
             �? i���t�?:            �X@"       #                    @M@�q�q�?             @������������������������       �                      @������������������������       �                     �?%       4                   �l@<����?8            �W@&       1       	          ����?(N:!���?'            �Q@'       *                   �X@     �?#             P@(       )                   �W@�����H�?
             2@������������������������       �        	             0@������������������������       �                      @+       0                    �?��<b�ƥ?             G@,       /                    �E@�g�y��?             ?@-       .                    @D@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     :@������������������������       �                     .@2       3                   �b@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     9@6       e                    �?���B���?�            �s@7       X                    �?�Y �K�?;            @X@8       =                    �?�A����?1            �T@9       :                    �M@�KM�]�?
             3@������������������������       �                     0@;       <                   `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?>       O                    �?�q�q�?'            �O@?       N       	          ����?��k=.��?            �G@@       C                   �e@���V��?            �F@A       B                   Pe@�q�q�?             @������������������������       �                     @������������������������       �                      @D       G                   `\@�ݜ�?            �C@E       F                   pb@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @H       I                   �c@(;L]n�?             >@������������������������       �        	             2@J       K                    b@�8��8��?             (@������������������������       �                     $@L       M                   8s@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @P       U                    �?      �?
             0@Q       R                   `k@�C��2(�?             &@������������������������       �                     @S       T                   n@      �?             @������������������������       �                     �?������������������������       �                     @V       W                    a@���Q��?             @������������������������       �                     @������������������������       �                      @Y       Z                    �?���Q��?
             .@������������������������       �                      @[       d                   �b@�	j*D�?             *@\       _       	          ����?      �?              @]       ^                    �?      �?             @������������������������       �                     �?������������������������       �                     @`       c                   �^@      �?             @a       b                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @f       w                     R@�?�|�?�            �k@g       h                    �J@ �Jj�G�?�            �k@������������������������       �        \            �b@i       v                   @g@����Q8�?-            �Q@j       q                   `d@hA� �?,            �Q@k       l       	            �?0�)AU��?"            �L@������������������������       �                    �I@m       p                    �?r�q��?             @n       o                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r       s                    c@8�Z$���?
             *@������������������������       �                     $@t       u                   0e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @y       �       
             �?�C�ӌ�?           p{@z       �                    �R@�&�TA�?�             w@{       �                   �c@�~Bo�?�            �v@|       �                   �`@0�b���?�            �t@}       �       	          `ff�?�"ZN��?^            �b@~       �                    �?>���a��?8            �V@       �                    �D@      �?              @������������������������       �                      @�       �       	             �?r�q��?             @������������������������       �                     @�       �                   (q@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          033�?�p ��?1            �T@�       �                    �?�>����?!             K@�       �                   �R@�IєX�?            �I@������������������������       �                     �?�       �                   �X@`2U0*��?             I@�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   (q@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �\@����?�?            �F@�       �                   �m@�IєX�?             1@�       �                    �J@      �?              @�       �                    �D@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     <@�       �                    @N@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    ]@����X�?             <@������������������������       �                     @�       �                   �_@���|���?             6@�       �                   �b@      �?              @�       �       
             �?      �?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    @d}h���?	             ,@�       �                    �N@�8��8��?             (@������������������������       �                     @�       �                   �_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �Z@XB���?&             M@�       �                   Pd@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   @\@@3����?#             K@�       �                   �o@�IєX�?
             1@������������������������       �                     &@�       �       	          ���@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                    �B@�       �                   0`@@>ZAɥ�?p            `g@�       �                   `Q@ 
�V�?R            �`@�       �                    �?�g�y��?             ?@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     <@������������������������       �        @            �Y@�       �                    �?�NW���?            �J@�       �                   �`@P�Lt�<�?             C@�       �                    �?�C��2(�?             &@������������������������       �                     @�       �       	             �?؇���X�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     ;@�       �                   �a@z�G�z�?	             .@�       �                   �n@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �q@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?���>4��?             <@�       �                    �?      �?              @������������������������       �                     @�       �                     I@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?���Q��?             4@�       �                   `l@X�<ݚ�?             2@������������������������       �                     @�       �                    �?�q�q�?	             (@������������������������       �                     @�       �                    @      �?              @�       �                   `\@z�G�z�?             @�       �                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �       	             @���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?\��_��?2            �Q@�       �                   `T@�8��8��?
             (@������������������������       �                     �?������������������������       �        	             &@�       �                    �?��Q:��?(            �M@�       �                    �?�GN�z�?             F@�       �                    �N@�n_Y�K�?             :@�       �                    @M@      �?             4@�       �                    `@X�Cc�?	             ,@������������������������       �                     @�       �                   0m@      �?             $@������������������������       �                     @�       �                   �e@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   Pa@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@�       �                    ]@z�G�z�?             .@������������������������       �                     �?�       �                   `f@؇���X�?             ,@������������������������       �                     (@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �x@     P�@     @t@     `c@     �E@     @]@      4@      (@      4@      @      4@      @      4@      @      4@       @              �?      4@      �?      @      �?       @      �?              �?       @              @              *@                      �?               @               @              @      7@     @Z@      *@      1@              &@      *@      @      (@      @      �?      @      �?                      @      &@              �?      @              @      �?              $@      V@       @      �?       @                      �?       @     �U@       @      O@      @     �N@       @      0@              0@       @              �?     �F@      �?      >@      �?      @              @      �?                      :@              .@      @      �?      @                      �?              9@     �q@      C@     @P@      @@     �M@      7@      1@       @      0@              �?       @               @      �?              E@      5@      C@      "@      C@      @      @       @      @                       @      A@      @      @      @      @                      @      =@      �?      2@              &@      �?      $@              �?      �?              �?      �?                       @      @      (@      �?      $@              @      �?      @      �?                      @      @       @      @                       @      @      "@       @              @      "@      @      @      �?      @      �?                      @      @      �?      �?      �?      �?                      �?       @                      @      k@      @      k@      @     �b@             �P@      @     �P@      @      L@      �?     �I@              @      �?      �?      �?              �?      �?              @              &@       @      $@              �?       @               @      �?                      �?               @      R@     �v@     �C@     �t@     �B@     `t@      8@     ps@      3@      `@      1@     @R@      @      @               @      @      �?      @               @      �?       @                      �?      (@     �Q@      @      I@      @      H@      �?               @      H@      �?      @               @      �?       @      �?                       @      �?      F@      �?      0@      �?      @      �?      @              @      �?                      @              "@              <@      �?       @      �?                       @       @      4@              @       @      ,@      @      @      @      @      @      �?              �?      @                       @       @              @      &@      �?      &@              @      �?      @              @      �?               @               @      L@      �?      @              @      �?              �?     �J@      �?      0@              &@      �?      @              @      �?                     �B@      @     �f@      �?     �`@      �?      >@      �?       @      �?                       @              <@             �Y@      @     �H@      �?     �B@      �?      $@              @      �?      @      �?       @      �?                       @              @              ;@      @      (@       @       @       @                       @      �?      $@              $@      �?              *@      .@      �?      @              @      �?      @      �?                      @      (@       @      $@       @      @              @       @              @      @      @      @      �?       @      �?              �?       @               @                      @       @               @      @       @                      @     �@@      C@      &@      �?              �?      &@              6@     �B@      $@      A@      $@      0@      $@      $@      @      "@              @      @      @              @      @      �?      @                      �?      @      �?      @                      �?              @              2@      (@      @              �?      (@       @      (@                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��{hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�<         �                    �?n[��L��?J           ��@       M       
             �?(�9�5�?.           0|@       D       	          pff�?4և����?�             u@       =                   �a@� ����?�             j@                           �?�iʫ{�?j            �c@                          �Z@b�2�tk�?             2@������������������������       �                     @                          �s@d}h���?
             ,@	       
                    �?      �?              @������������������������       �                      @                           �?      �?             @������������������������       �                      @              	          433�?      �?             @������������������������       �                      @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       :                   �e@Tri����?^            �a@       !                    @L@�θV�?\            @a@              
             �?Х-��ٹ?1            �R@������������������������       �                     @                           l@ >�֕�?,            �Q@������������������������       �                    �D@                            �?\-��p�?             =@                           \@ �Cc}�?             <@������������������������       �                     �?                          ``@�>����?             ;@������������������������       �                     ,@                           @H@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     �?"       +                    �?��d��?+            �O@#       &       
             �?�z�G��?             4@$       %                    @P@      �?             @������������������������       �                      @������������������������       �                      @'       *                   �q@      �?             0@(       )                   0a@؇���X�?             ,@������������������������       �        
             (@������������������������       �                      @������������������������       �                      @,       5       	          `ff�?�ʈD��?            �E@-       4                    [@�IєX�?             A@.       /                   @_@r�q��?             (@������������������������       �                     @0       1                    �N@�q�q�?             @������������������������       �                      @2       3                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     6@6       7                   �^@�<ݚ�?             "@������������������������       �                     @8       9                    @M@�q�q�?             @������������������������       �                      @������������������������       �                     �?;       <                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @>       C                    �?`2U0*��?"             I@?       B                    �M@z�G�z�?             $@@       A                   Pt@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     D@E       L                    \@����}��?S            �_@F       K                   �_@������?             B@G       H                   �o@r�q��?             @������������������������       �                     @I       J                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     >@������������������������       �        ;            �V@N       s       	          ����?�2��P��?O            �\@O       Z                   �b@���"͏�?4            �R@P       W                    �?�q��/��?             G@Q       R                    X@@-�_ .�?            �B@������������������������       �                     �?S       V                    �?������?             B@T       U                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                    �@@X       Y                   �^@�q�q�?             "@������������������������       �                     @������������������������       �                     @[       \                   �e@���>4��?             <@������������������������       �                     @]       h                   8q@      �?             8@^       g                    �L@z�G�z�?
             .@_       f                   �l@؇���X�?	             ,@`       e                    �?�<ݚ�?             "@a       b                   @i@����X�?             @������������������������       �                     �?c       d                   �a@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?i       p                    �?�q�q�?             "@j       o                   0w@����X�?             @k       n                    �?r�q��?             @l       m                    d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     �?q       r                   c@      �?              @������������������������       �                     �?������������������������       �                     �?t       w                    �?� ��1�?            �D@u       v                    `@      �?             @������������������������       �                      @������������������������       �                      @x       {                    �?�MI8d�?            �B@y       z                   c@      �?	             (@������������������������       �                     "@������������������������       �                     @|       }       	          033�?H%u��?             9@������������������������       �                     ,@~              	          ����?���!pc�?             &@������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     @�       �                   �_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    I@�zFn��?           0}@�       �                   �e@�<ݚ�?            �F@�       �       	          033�?&^�)b�?            �E@�       �                   �b@l��
I��?             ;@�       �       
             �?�+e�X�?             9@������������������������       �                      @�       �       
             �?�㙢�c�?             7@�       �                   �^@�}�+r��?             3@�       �                   �Z@�����H�?             "@�       �                    @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@������������������������       �                      @�       �                    �K@PB�~�?�            `z@�       �       	          ����?������?�            �q@�       �                   �z@Du9iH��?�            �j@�       �                    @@�S�1�?             j@�       �       	          ����?` A�c̭?y             i@�       �                   h@��8����?t             h@�       �                    �? ������?r            �g@�       �                    �?`��>�ϗ?g            @e@�       �                   �a@ A��� �?b            @d@�       �                     B@�Ń��̧?             E@������������������������       �                     �?������������������������       �                    �D@������������������������       �        E             ^@�       �                   �q@      �?              @������������������������       �                     @������������������������       �                     �?�       �                   �m@�}�+r��?             3@������������������������       �                     "@�       �       
             �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                   �h@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    a@      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             "@������������������������       �                     @�       �       
             �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?@i��M��?*            @P@�       �                    b@      �?             8@�       �                    �?���7�?             6@������������������������       �                     0@�       �                   �\@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       	          ����?�>$�*��?            �D@�       �                   �q@z�G�z�?             $@�       �                   �b@�����H�?             "@������������������������       �                     @�       �                   @c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �       
             �?�4�����?             ?@�       �       
             �?\X��t�?             7@������������������������       �                     @�       �                    �?      �?             4@������������������������       �                     @�       �                     F@�q�q�?             .@������������������������       �                     @�       �                    n@�C��2(�?	             &@������������������������       �                     @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�                          �?L�];�?T            �a@�       �                    q@��ɜ|��?>            �Z@�       �                    `@z\�3�?,            �S@������������������������       �                     ,@�       �       	          033@�	j*D�?$            @P@�       �                   �X@ {��e�?            �J@������������������������       �                     @�       �                    @M@�J�4�?             I@�       �                    �?�	j*D�?             *@������������������������       �                     @�       �                    �L@ףp=
�?             $@������������������������       �                      @�       �                    m@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   0c@������?            �B@�       �                   �k@8�Z$���?             :@�       �       
             �?      �?
             0@������������������������       �                     �?�       �       	          ����?z�G�z�?	             .@�       �                    �?և���X�?             @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     &@�       �       
             �?      �?             (@������������������������       �                     @������������������������       �                     "@�             	          ����?և���X�?             <@�                          @D�n�3�?             3@�       �                    �?     ��?             0@�       �                    �?r�q��?	             (@������������������������       �                     @�       �                   @c@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   @a@      �?             @������������������������       �                      @                         �u@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        pz@�����H�?             "@������������������������       �                      @������������������������       �                     �?            
             �?">�֕�?            �A@      	                   @M@��a�n`�?             ?@������������������������       �                     @
                        �\@ �o_��?             9@������������������������       �                     @                         �M@"pc�
�?             6@������������������������       �                     @                         �?�}�+r��?             3@������������������������       �                     *@                          O@r�q��?             @                        0b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�BP       �z@     �~@     �W@     Pv@      >@      s@      =@     �f@      ;@     �`@      &@      @              @      &@      @      @      @       @              @      @       @              �?      @               @      �?      �?              �?      �?              @              0@     @_@      ,@      _@      @     �Q@              @      @     �P@             �D@      @      9@      @      9@      �?               @      9@              ,@       @      &@              &@       @              �?              $@     �J@      @      ,@       @       @       @                       @      @      (@       @      (@              (@       @               @              @     �C@       @      @@       @      $@              @       @      @               @       @       @       @                       @              6@       @      @              @       @      �?       @                      �?       @      �?              �?       @               @      H@       @       @       @      �?              �?       @                      @              D@      �?     �_@      �?     �A@      �?      @              @      �?      �?              �?      �?                      >@             �V@      P@     �I@      L@      2@     �D@      @     �A@       @              �?     �A@      �?       @      �?       @                      �?     �@@              @      @              @      @              .@      *@              @      .@      "@      (@      @      (@       @      @       @      @       @              �?      @      �?      @                      �?       @              @                      �?      @      @       @      @      �?      @      �?      @      �?                      @               @      �?              �?      �?              �?      �?               @     �@@       @       @               @       @              @      ?@      @      "@              "@      @              @      6@              ,@      @       @       @              �?       @              @      �?      @              @      �?              u@     ``@      $@     �A@       @     �A@       @      3@      @      3@       @              @      3@      �?      2@      �?       @      �?       @               @      �?                      @              $@      @      �?      @                      �?       @                      0@       @             `t@      X@     �n@      B@      i@      .@      i@      "@     @h@      @     `g@      @     @g@      @      e@       @      d@      �?     �D@      �?              �?     �D@              ^@              @      �?      @                      �?      2@      �?      "@              "@      �?              �?      "@              �?       @               @      �?              @      �?      @                      �?      @      @      @               @      @              @       @                      @      F@      5@      5@      @      5@      �?      0@              @      �?              �?      @                       @      7@      2@       @       @      �?       @              @      �?       @      �?                       @      �?              5@      $@      *@      $@      @              $@      $@      @              @      $@      @              �?      $@              @      �?      @      �?                      @       @             �T@      N@     �Q@      B@     �M@      4@      ,@             �F@      4@      E@      &@              @      E@       @      "@      @              @      "@      �?       @              �?      �?              �?      �?             �@@      @      6@      @      (@      @              �?      (@      @      @      @      @              �?      @              @      �?               @              $@              &@              @      "@      @                      "@      (@      0@      &@       @      &@      @      $@       @      @              @       @      @                       @      �?      @               @      �?      �?              �?      �?                      @      �?       @               @      �?              &@      8@      @      8@              @      @      2@      @              @      2@      @              �?      2@              *@      �?      @      �?       @               @      �?                      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�WtNhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�6         t       	          ����?��J�0�?J           ��@       )       
             �?�!�����?6           �}@                            �?f1r��g�?m            �c@       	                   �`@�]F���?H            �Z@                          �X@ qP��B�?            �E@                           X@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                    �A@
                           �?     8�?-             P@                           �?@�0�!��?             A@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?              	          833�?��� ��?             ?@������������������������       �                     ;@������������������������       �                     @                          @j@      �?             >@������������������������       �                     @              	          ����?�LQ�1	�?             7@������������������������       �        	             "@              	          833�?և���X�?	             ,@                          �b@r�q��?             @������������������������       �                     @������������������������       �                     �?                          �l@      �?              @������������������������       �                     �?                           �K@����X�?             @              	          ����?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @!       "                    �? ��WV�?%             J@������������������������       �                     @#       $       	          833�?`�q�0ܴ?!            �G@������������������������       �                     C@%       (                   �[@�<ݚ�?             "@&       '                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @*       =                    �?أp=
��?�             t@+       4                   Hq@p�ݯ��?             �L@,       -                   0c@���?            �D@������������������������       �        	             .@.       3                   �[@�n_Y�K�?             :@/       0                    �H@r�q��?             (@������������������������       �                     @1       2                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             ,@5       :                    �?     ��?
             0@6       9                    d@�C��2(�?             &@7       8                   �c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @;       <                   �s@z�G�z�?             @������������������������       �                     @������������������������       �                     �?>       A                   �X@��.���?�            pp@?       @                    �I@      �?             $@������������������������       �                     @������������������������       �                     @B       [                    �?<��ٵ�?�            �o@C       V                    b@L=�m��?&            �N@D       K                   `]@؇���X�?"             L@E       J                   `\@�n_Y�K�?
             *@F       I                   �b@���!pc�?             &@G       H                   `X@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @L       O                   @E@Du9iH��?            �E@M       N                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @P       Q                    @M@�(\����?             D@������������������������       �                     B@R       U       	          ����?      �?             @S       T                    @N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @W       Z                   �d@���Q��?             @X       Y                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?\       m                    �O@      �?}             h@]       h       	            �?�ګ���?u            `f@^       g       	          ����?@c����?p            @e@_       `                    �?��ꤘ�?e             c@������������������������       �        ?            �X@a       f                   @[@@3����?&             K@b       e                    @r�q��?             @c       d                    c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        !             H@������������������������       �                     1@i       l       	          pff�?�����H�?             "@j       k                   @k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @n       s                   @t@�	j*D�?             *@o       p                    �?ףp=
�?             $@������������������������       �                     @q       r                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @u       �                    �?�C*�%��?           p{@v       �       	          `ff@؀�:M�?.            �R@w       �       
             �?�q�q�?*            @Q@x       �                   �b@X��ʑ��?            �E@y       �                   w@      �?             @@z       }                    @K@
;&����?             7@{       |                    @I@z�G�z�?             @������������������������       �                     �?������������������������       �                     @~       �                    @X�<ݚ�?             2@       �                    `@j���� �?             1@�       �                    �?�q�q�?	             (@�       �                   �`@���|���?             &@�       �                    �?؇���X�?             @������������������������       �                     @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                    �?�C��2(�?             &@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   ``@$�q-�?             :@�       �                   @]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     7@������������������������       �                     @�       �       	          ����?�d�QDn�?�            �v@�       �                   @h@��X���?/            @Q@�       �                    c@ 7���B�?             ;@������������������������       �                     9@�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �e@����X�?             E@�       �       
             �?      �?             D@�       �                    �?�>4և��?             <@�       �                   @k@ȵHPS!�?             :@�       �                    @K@      �?             @�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     4@������������������������       �                      @�       �                    �?�q�q�?	             (@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �c@����?�            �r@�       �                    @؝�x�O�?�            �p@�       �                   �Z@     ��?�             p@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �_@�nkK�?�            �o@�       �       
             �?���}<S�?'            @Q@�       �                    �?��S�ۿ?"             N@�       �                    @P@�&=�w��?            �J@�       �       	             �?@��8��?             H@�       �                     F@�nkK�?             7@�       �                   �\@      �?             @������������������������       �                     �?�       �                   c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             3@������������������������       �                     9@�       �                   �\@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �^@����X�?             @������������������������       �                     @������������������������       �                      @�       �                    �H@�<ݚ�?             "@������������������������       �                     �?�       �                    ]@      �?              @������������������������       �                      @�       �                   `U@r�q��?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       
             �?�˫���?t             g@�       �                     E@�Sa��?k            �d@�       �                    b@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    c@�dJ�Ҙ?h            `d@������������������������       �        c            �b@�       �                    �?؇���X�?             ,@������������������������       �                     @�       �                   pc@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�       �                   �a@�t����?	             1@�       �                   c@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@�       �       
             �?�	j*D�?             *@�       �       	          `ff�?"pc�
�?             &@������������������������       �                     @�       �       
             �?����X�?             @������������������������       �                     �?�       �                    ^@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?�q�q�?             ;@�       �                    ]@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �E@��.k���?
             1@������������������������       �                     @�       �                    �J@X�Cc�?             ,@������������������������       �                     @�       �                    b@�eP*L��?             &@�       �                   �d@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�        x@     ��@     �r@     @f@      8@     �`@      6@     @U@      �?      E@      �?      @              @      �?                     �A@      5@     �E@      @      <@       @      �?       @                      �?      @      ;@              ;@      @              .@      .@      @               @      .@              "@       @      @      @      �?      @                      �?      @      @      �?               @      @       @       @       @                       @              @       @      I@              @       @     �F@              C@       @      @       @      �?       @                      �?              @     Pq@     �E@      B@      5@      ?@      $@      .@              0@      $@       @      $@              @       @      @              @       @              ,@              @      &@      �?      $@      �?      @              @      �?                      @      @      �?      @                      �?      n@      6@      @      @      @                      @     �m@      1@      I@      &@      H@       @       @      @       @      @       @      �?              �?       @                       @               @      D@      @      �?       @      �?                       @     �C@      �?      B@              @      �?      �?      �?              �?      �?               @               @      @      �?      @              @      �?              �?             @g@      @      f@       @      e@      �?      c@      �?     �X@             �J@      �?      @      �?      @      �?              �?      @               @              H@              1@               @      �?      �?      �?      �?                      �?      @              "@      @      "@      �?      @               @      �?       @                      �?              @     @U@      v@      G@      <@      G@      7@      6@      5@      (@      4@      (@      &@      @      �?              �?      @               @      $@      @      $@      @      @      @      @      @      �?      @              �?      �?              �?      �?              �?      @              @      �?                      �?              @      �?                      "@      $@      �?      �?      �?      �?                      �?      "@              8@       @      �?       @      �?                       @      7@                      @     �C@     `t@      *@      L@      �?      :@              9@      �?      �?              �?      �?              (@      >@      $@      >@      @      7@      @      7@      @      @      �?      @               @      �?      �?      �?                      �?       @                      4@       @              @      @      �?      @              @      �?              @               @              :@     �p@      1@     �o@      *@     `n@       @      �?       @                      �?      &@     @n@      @     �O@      @      L@       @     �I@      �?     �G@      �?      6@      �?      @              �?      �?       @      �?                       @              3@              9@      �?      @      �?                      @       @      @              @       @               @      @      �?              �?      @               @      �?      @      �?      @      �?                      @               @      @     `f@      @     �d@      �?      @              @      �?               @      d@             �b@       @      (@              @       @      @       @                      @       @      .@       @      @              @       @                      $@      @      "@       @      "@              @       @      @      �?              �?      @      �?                      @       @              "@      2@      �?      "@      �?                      "@       @      "@      @              @      "@              @      @      @       @      @       @                      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��8hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK酔h~�B�2         T       	          ����?X�<ݚ�??           ��@       !       
             �?���m��?           �{@              	          ����?��\���?U            @`@                          �b@�8��8��?J             [@       
                   `\@ ��N8�?8             U@                           T@�C��2(�?             &@������������������������       �                      @       	                   `f@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        1            @R@                           �?�q�q�?             8@                          `]@��.k���?             1@������������������������       �                     @                           @C@�n_Y�K�?
             *@������������������������       �                      @                           �?���!pc�?             &@                          �i@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @                          ``@���|���?             6@                          �c@z�G�z�?             .@������������������������       �                     $@                           �?���Q��?             @������������������������       �                      @������������������������       �                     @                            �?����X�?             @                            F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @"       =                    �L@P5�޷�?�            �s@#       $                    �?`Jj��?�             o@������������������������       �        ,            �Q@%       6                    �?�����?j             f@&       '                    X@��[�8��?            �I@������������������������       �                     @(       )                    �A@r�q��?             H@������������������������       �                     �?*       -                    P@��0{9�?            �G@+       ,                   p`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @.       5                    �?@4և���?             E@/       0                   �e@l��\��?             A@������������������������       �                     =@1       4                   �`@���Q��?             @2       3                   �f@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @7       8                    @G@ ,V�ނ�?K            �_@������������������������       �        (             P@9       <                    �G@6uH���?#             O@:       ;                   @[@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      K@>       K                   �b@���!pc�?%            �P@?       J                   �j@r�q��?             E@@       E                    �?j���� �?             1@A       D       	            �?�q�q�?             "@B       C                   �a@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @F       I       	          ����?      �?              @G       H                    ^@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     9@L       S                    �?r�q��?             8@M       R                   �e@ҳ�wY;�?
             1@N       O                    �?������?	             .@������������������������       �                     "@P       Q                    @N@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @U       �                   �b@L�Sg��?/           �}@V       �                    �?,���i�?�            w@W       X                   �U@t-+��?�            pr@������������������������       �                      @Y       �                    �R@��Xb�?�            Pr@Z       q                   `_@�L�A�?�             r@[       h       	          ����?0���ަ?l            �e@\       a                    �?0G���ջ?              J@]       `                    �?      �?             @^       _                    �N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?b       c                    �?@��8��?             H@������������������������       �                    �C@d       e                    �?�����H�?             "@������������������������       �                     �?f       g                   �X@      �?              @������������������������       �                     �?������������������������       �                     @i       j       	          `ff@ �|ك�?L            �^@������������������������       �        B            �Z@k       l                    �?�IєX�?
             1@������������������������       �                     &@m       p       	          ���	@r�q��?             @n       o                     M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @r                          �b@d����?M            �\@s       ~                    �L@Pq�����?9            @U@t       y                   �\@HP�s��?!             I@u       x       	          ����?      �?              @v       w                   @Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @z       {                   r@�Ń��̧?             E@������������������������       �                     A@|       }                    �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                    �A@�       �       
             �?�z�G��?             >@�       �                    �?���B���?             :@�       �       
             �?���|���?             &@������������������������       �                      @�       �                    �?X�<ݚ�?             "@������������������������       �                      @�       �                   `c@և���X�?             @������������������������       �                     @�       �       	          ����?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?��S�ۿ?             .@�       �                    `@r�q��?             @�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     @�       �                   n@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?4�B��?0            �R@�       �                    \@���Q��?"            �K@�       �                   @_@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��H�}�?             I@�       �                    �K@؇���X�?             @������������������������       �                     @�       �                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �e@^����?            �E@�       �                   �_@���?            �D@�       �                    @�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�       �                   P`@8^s]e�?             =@�       �       	          ����?�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �       
             �?R���Q�?             4@������������������������       �                      @�       �                    @M@�X�<ݺ?             2@������������������������       �                     $@�       �                     P@      �?              @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   @_@�KM�]�?             3@�       �                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �R@�IєX�?             1@������������������������       �                     0@������������������������       �                     �?�       �                   Pc@և���X�?C            @Z@�       �                   �w@�IєX�?             1@������������������������       �        
             0@������������������������       �                     �?�       �       
             �?      �?8             V@�       �                    �?N{�T6�?"            �K@�       �                   �q@�p ��?            �D@�       �                   g@����e��?            �@@�       �       	             @f���M�?             ?@�       �       	          ����?      �?             6@�       �                    �?ҳ�wY;�?             1@�       �                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   0`@����X�?             ,@�       �                    @E@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                    @K@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     "@������������������������       �                      @������������������������       �                      @������������������������       �                     ,@�       �       	          033@:ɨ��?            �@@�       �                     M@r֛w���?             ?@�       �                    �F@r�q��?             8@������������������������       �                      @�       �                   �d@      �?
             0@�       �                    �?�C��2(�?             &@������������������������       �                      @�       �                    �?�q�q�?             @�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   pg@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       	          033�?և���X�?             @�       �                   �t@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�t�b�$     h�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@     �r@     �a@      7@     �Z@      "@     �X@      �?     �T@      �?      $@               @      �?       @      �?                       @             @R@       @      0@       @      "@              @       @      @               @       @      @       @      �?              �?       @                       @              @      ,@       @      (@      @      $@               @      @       @                      @       @      @       @      �?              �?       @                      @     �q@      A@      m@      0@     �Q@              d@      0@      D@      &@              @      D@       @              �?      D@      @      �?      @      �?                      @     �C@      @      ?@      @      =@               @      @       @      �?              �?       @                       @       @             @^@      @      P@             �L@      @      @      @              @      @              K@              H@      2@     �A@      @      $@      @      @      @      �?      @              @      �?               @              @      �?      @      �?      @                      �?      @              9@              *@      &@      @      &@      @      &@              "@      @       @               @      @               @              @             @Z@     w@     �F@     @t@      5@      q@       @              3@      q@      1@     q@      @     `e@      @     �H@       @       @      �?       @      �?                       @      �?              �?     �G@             �C@      �?       @              �?      �?      @      �?                      @      �?     �^@             �Z@      �?      0@              &@      �?      @      �?      �?      �?                      �?              @      *@     �Y@      @     @T@      @      G@      @      @      @      �?              �?      @                      @      �?     �D@              A@      �?      @      �?                      @             �A@      "@      5@      @      5@      @      @               @      @      @               @      @      @      @              �?      @      �?                      @      �?      ,@      �?      @      �?      �?      �?                      �?              @              "@      @               @      �?              �?       @              8@      I@      6@     �@@      @      �?      @                      �?      2@      @@      @      �?      @               @      �?              �?       @              (@      ?@      $@      ?@      �?      &@              &@      �?              "@      4@      @      @              @      @              @      1@       @              �?      1@              $@      �?      @      �?      �?              �?      �?                      @       @               @      1@      �?      �?              �?      �?              �?      0@              0@      �?              N@     �F@      0@      �?      0@                      �?      F@      F@      5@      A@      5@      4@      *@      4@      &@      4@      &@      &@      @      &@       @      �?              �?       @              @      $@      �?       @      �?                       @      @       @               @      @              @                      "@       @               @                      ,@      7@      $@      7@       @      4@      @       @              (@      @      $@      �?       @               @      �?      �?      �?      �?                      �?      �?               @      @       @                      @      @      @      �?      @              @      �?               @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��(hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�Bx=         t                   �`@�	����?C           ��@       '       	          ����?���G�?           {@              
             �? �q(���?c            �c@                           �?��(\���?3             T@                          �_@      �?              H@                           @L@���N8�?             E@                           �?�KM�]�?             3@       	                   0l@$�q-�?
             *@������������������������       �                      @
                           \@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                          �X@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     7@                           _@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @@              	             �$��$�L�?0            �S@������������������������       �                      @       $                   �S@�S(��d�?/            @S@                           @I@�q�q�?             (@������������������������       �                      @                           �?      �?             $@                           �?z�G�z�?             @                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?        !                   �a@z�G�z�?             @������������������������       �                      @"       #                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?%       &                    @ ����?'            @P@������������������������       �        &             P@������������������������       �                     �?(       A                    �?��)��g�?�             q@)       *                   @W@��6}��?%            �N@������������������������       �                     @+       6       	          pff�?����X�?!             L@,       -                    �?      �?             4@������������������������       �                     @.       /                   �]@�θ�?             *@������������������������       �                     @0       1                   @_@      �?             @������������������������       �                      @2       3                    b@      �?             @������������������������       �                      @4       5       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?7       >                   �r@r�q��?             B@8       =                    �?      �?             @@9       <       	          ����?���y4F�?             3@:       ;       	          033�?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     $@������������������������       �                     *@?       @                     J@      �?             @������������������������       �                      @������������������������       �                      @B       I                   �[@�����?�            �j@C       H                   �[@`����֜?0            �Q@D       G                   �Y@؇���X�?             @E       F                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        +            �O@J       U                    \@�1�hP	�?Y            �a@K       L                   Pn@�q�q�?	             .@������������������������       �                     @M       N       	             �?�eP*L��?             &@������������������������       �                     �?O       T                    �?      �?             $@P       Q                     M@      �?              @������������������������       �                     @R       S                   �q@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @V       q                    @     p�?P             `@W       j       
             �?H�̱���?N            @_@X       ]                    @H@����w�?F            @[@Y       \       	          ����?�KM�]�?             3@Z       [                   `\@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     .@^       a                    �?����?�?;            �V@_       `       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @b       i                   P`@���E�?8            �U@c       d                    @M@ 7���B�?             ;@������������������������       �                     5@e       f                   �_@r�q��?             @������������������������       �                     @g       h                   �r@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        (             N@k       l                   �_@      �?             0@������������������������       �                     @m       p                   �r@X�<ݚ�?             "@n       o                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @r       s                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?u       �                    �K@`��t��?2           P~@v       �                    �?hBW�=��?�            `u@w       �       	          hff�?�Ƀ aA�?L            �]@x                          �b@�6����?,            @R@y       ~                    �G@�S����?             3@z       {                   0a@      �?             (@������������������������       �                      @|       }                   �a@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @�       �                   `@���3L�?             K@�       �                   �f@V�a�� �?             =@�       �                    \@PN��T'�?             ;@�       �                     H@������?             .@�       �                    �E@8�Z$���?             *@�       �                    �?����X�?             @������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                     �?�       �                    �D@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     (@������������������������       �                      @�       �                   pf@`�Q��?             9@�       �                    �?�<ݚ�?             2@�       �       
             �?��S�ۿ?             .@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                     @�       �                   @b@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �e@��Hg���?             �F@�       �                   �\@d}h���?             E@�       �                   �b@���Q��?             $@������������������������       �                     @������������������������       �                     @�       �                    �J@     ��?             @@�       �                   �g@`2U0*��?             9@�       �                   �e@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     4@�       �       
             �?����X�?             @������������������������       �                     @������������������������       �                      @�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       
             �?     ��?�             l@�       �                    �?�q�q�?!             H@�       �                   �b@$�q-�?             *@������������������������       �        
             (@������������������������       �                     �?�       �                    �?�xGZ���?            �A@�       �                   g@l��
I��?             ;@�       �                    �E@�+e�X�?             9@�       �                   @_@և���X�?             @�       �                   `e@�q�q�?             @�       �                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   0f@r�q��?             2@�       �                    �?�t����?
             1@������������������������       �                     �?�       �                    b@      �?	             0@�       �       	          ����?z�G�z�?             @�       �                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �? J���#�?e             f@�       �                   �p@�nkK�?             7@������������������������       �        	             ,@�       �                   �g@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �        V             c@�                          �?��O�A�?`            �a@�       �                    �?�o;����?<            �S@�       �                   �a@������?*             L@������������������������       �                     (@�       �                    �?~�4_�g�?#             F@�       �       	          ����?��H�}�?             9@�       �                   �q@     ��?             0@�       �                   �m@�z�G��?             $@�       �                   pd@���Q��?             @�       �                    @L@�q�q�?             @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     @�       �                   0r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@�       �                    @N@�S����?             3@�       �                    @L@�q�q�?             "@�       �                    �?z�G�z�?             @�       �                   8p@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �       
             �?      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                    �?8����?             7@������������������������       �                     "@�       �                    @O@      �?             ,@�       �                    @�q�q�?	             "@�       �                   @a@����X�?             @������������������������       �                     @�       �       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?                         �d@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                        �^@     ��?$             P@            
             �?��S���?             .@������������������������       �                     @                        �]@�q�q�?             (@      
                   �O@X�<ݚ�?             "@      	                   �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @                        `f@��<D�m�?            �H@            
             �?�(\����?             D@������������������������       �                    �@@                         �?؇���X�?             @������������������������       �                     @������������������������       �                     �?                         c@�<ݚ�?             "@            	          ����?      �?              @                        �g@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KMKK��h_�B�        z@     `@     @[@     @t@     @S@     �T@      @     �R@      @      E@       @      D@       @      1@      �?      (@               @      �?      @      �?                      @      �?      @      �?                      @              7@      @       @               @      @                      @@     �Q@       @               @     �Q@      @      @      @       @              @      @      @      �?      @      �?              �?      @              �?              �?      @               @      �?       @               @      �?              P@      �?      P@                      �?      @@     @n@      0@     �F@              @      0@      D@      $@      $@      @              @      $@              @      @      @       @              �?      @               @      �?      �?              �?      �?              @      >@      @      <@      @      .@      @      @              @      @                      $@              *@       @       @               @       @              0@     �h@      �?     @Q@      �?      @      �?      �?              �?      �?                      @             �O@      .@      `@      @      $@              @      @      @              �?      @      @      @      @      @               @      @              @       @                       @      $@     �]@       @     @]@      @     @Z@       @      1@       @       @               @       @                      .@       @      V@      �?       @      �?                       @      �?     �U@      �?      :@              5@      �?      @              @      �?       @               @      �?                      N@      @      (@              @      @      @      @      �?              �?      @                      @       @      �?       @                      �?     0s@     @f@     �o@     @V@      I@      Q@     �C@      A@      0@      @      "@      @               @      "@      �?      "@                      �?      @              7@      ?@      @      7@      @      7@      @      &@       @      &@       @      @               @       @      @              �?       @       @               @       @                      @       @                      (@       @              1@       @      ,@      @      ,@      �?      @      �?      @                      �?      &@                      @      @      @      @                      @      &@      A@      "@     �@@      @      @      @                      @      @      =@      �?      8@      �?      @              @      �?                      4@       @      @              @       @               @      �?              �?       @             `i@      5@      <@      4@      (@      �?      (@                      �?      0@      3@       @      3@      @      3@      @      @       @      @       @      �?              �?       @                      @      �?              @      .@       @      .@      �?              �?      .@      �?      @      �?      �?      �?                      �?              @              &@      �?               @               @             �e@      �?      6@      �?      ,@               @      �?       @                      �?      c@              K@     @V@      F@     �A@     �B@      3@      (@              9@      3@      "@      0@      "@      @      @      @       @      @       @      �?      �?              �?      �?              �?      �?                       @      @               @      @              @       @      �?              �?       @                      "@      0@      @      @      @      @      �?      @      �?      @                      �?      �?               @       @      �?              �?       @              �?      �?      �?      �?                      �?      $@              @      0@              "@      @      @      @      @       @      @              @       @      �?              �?       @              �?      �?              �?      �?              @      �?      @                      �?      $@      K@      @       @              @      @      @      @      @       @      @              @       @               @              @              @      G@      �?     �C@             �@@      �?      @              @      �?               @      @      �?      @      �?      @      �?                      @              @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJE�FhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B�4         �       
             �?�5��?N           ��@       Q                    �?�5�ط^�?\           ��@                           @G@�)���Y�?�            �x@       	                    �?&�a2o��?$            @Q@                          �a@"pc�
�?             &@                           �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     �?
                          �e@�y��*�?             M@                           @D@,�+�C�?            �K@������������������������       �                     9@                           �?�r����?             >@                          pb@�����H�?             ;@������������������������       �                     6@                           `@���Q��?             @������������������������       �                     @������������������������       �                      @                          �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @              	          833�?>iFa��?�            0t@������������������������       �        &            �N@       H                    �?0�v���?�            `p@       !       	          pff�?�wV����?r            �e@                          �X@���!pc�?             &@������������������������       �                      @              	          ����?�����H�?             "@������������������������       �                     @                            �L@      �?             @������������������������       �                     �?������������������������       �                     @"       ;                    �?����?j            �d@#       $                   �V@H�Swe�?S            @_@������������������������       �                     �?%       &                   @^@`�c�г?R             _@������������������������       �        &            �O@'       2                    �?85�}C�?,            �N@(       1                   �a@z�G�z�?             .@)       .                   �^@�q�q�?             "@*       +       	             �?�q�q�?             @������������������������       �                     �?,       -                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?/       0                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @3       :                   pi@�nkK�?              G@4       5                    ^@z�G�z�?             $@������������������������       �                     �?6       7                   �V@�����H�?             "@������������������������       �                     @8       9                   �g@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     B@<       G                   �p@�ݜ�?            �C@=       F                   @^@z�G�z�?             9@>       ?       
             �?�q�q�?             (@������������������������       �                     �?@       E       	             @���|���?             &@A       B                   �_@���Q��?             $@������������������������       �                      @C       D                   �X@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                     ,@I       P                    �?���E�?4            �U@J       K                    �?@��8��?              H@������������������������       �                     $@L       O       
             �?P�Lt�<�?             C@M       N                   �a@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @@������������������������       �                    �C@R       �                    �?�!���?l            @e@S       ^                    �?���b���?H            �\@T       W                   ph@      �?             4@U       V                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?X       Y                   pm@@�0�!��?             1@������������������������       �                     @Z       ]       	             �?�z�G��?             $@[       \                   �p@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @_       z                   a@z�J�?9            �W@`       o                   Pd@~|z����?#            �J@a       j       	          ����?���!pc�?            �@@b       c                   `X@D�n�3�?             3@������������������������       �                     @d       g                    �?     ��?             0@e       f                     C@z�G�z�?             @������������������������       �                     �?������������������������       �                     @h       i       	          ����?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?k       l                    �?@4և���?             ,@������������������������       �        	             (@m       n                    @      �?              @������������������������       �                     �?������������������������       �                     �?p       q                   @W@z�G�z�?             4@������������������������       �                      @r       y                    �L@�����H�?             2@s       t                   �e@�IєX�?
             1@������������������������       �                      @u       x       	          ����?�����H�?             "@v       w                    ]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?{       �                    �?�p ��?            �D@|       }       
             �?���Q��?
             .@������������������������       �                     @~       �                   �a@      �?             (@       �                    @�q�q�?             @������������������������       �                     �?�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     O@�����H�?             "@������������������������       �                     @�       �                   pk@      �?             @������������������������       �                      @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     :@�       �                   �[@�X�C�?$             L@�       �       	          @33�?      �?              @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     @�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `c@      �?             H@�       �       	          ����?`�q�0ܴ?            �G@�       �                   �`@ףp=
�?             4@������������������������       �        
             1@�       �                   pa@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ;@������������������������       �                     �?�       �                   @E@~�dis��?�            @v@�       �                    �?��[�p�?            �G@�       �                    �?�\��N��?             3@�       �                     F@z�G�z�?             $@�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     @�       �       	          ����?�<ݚ�?             "@�       �                    �?���Q��?             @�       �                    \@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     <@�       �                    �?\�t��Y�?�            Ps@�       �                   �g@�iyw	
�?�            �p@�       �                    @L@�{��?�            �p@�       �                   �[@�#w
:��?�            �i@�       �                    �?@4և���?             <@�       �                    �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     5@�       �                    �?�O"9��?{             f@�       �                    �I@г�wY;�?             A@������������������������       �                     :@�       �                   �_@      �?              @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        a            �a@�       �       	             @��a�n`�?.             O@�       �       	          833�?��f/w�?-            �N@�       �                    b@�E��ӭ�?             B@�       �                    �?д>��C�?             =@�       �                    �?�E��ӭ�?             2@�       �                    �?      �?             @�       �                   �p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    c@؇���X�?
             ,@������������������������       �                     $@�       �                    �?      �?             @�       �                   f@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     &@�       �                    ^@����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?H%u��?             9@������������������������       �                     @�       �                     M@r�q��?             2@������������������������       �                     �?�       �                   �c@�t����?             1@�       �                    �?      �?             0@�       �                   �n@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �?�>$�*��?            �D@�       �                    �?      �?             8@�       �                    �?�d�����?
             3@�       �                    �?�q�q�?             (@������������������������       �                     @�       �       	          ����?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �`@z�G�z�?             @������������������������       �                     @�       �                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     1@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B       `w@      �@     �V@     p}@      B@     @v@      0@     �J@      "@       @      "@      �?      "@                      �?              �?      @     �I@      @     �I@              9@      @      :@      @      8@              6@      @       @      @                       @      �?       @               @      �?              @              4@     �r@             �N@      4@     @n@      3@     �c@       @      @               @       @      �?      @              @      �?              �?      @              &@      c@      @     �]@      �?              @     �]@             �O@      @      L@      @      (@      @      @       @      �?      �?              �?      �?              �?      �?              �?      @      �?                      @              @       @      F@       @       @      �?              �?       @              @      �?      @      �?                      @              B@      @      A@      @      4@      @      @      �?              @      @      @      @       @               @      @       @                      @              �?              *@              ,@      �?     �U@      �?     �G@              $@      �?     �B@      �?      @              @      �?                      @@             �C@     �K@     �\@      G@      Q@      .@      @      �?       @               @      �?              ,@      @      @              @      @      @      @              @      @              @              ?@     �O@      9@      <@      "@      8@       @      &@      @              @      &@      @      �?              �?      @              �?      $@              $@      �?              �?      *@              (@      �?      �?      �?                      �?      0@      @               @      0@       @      0@      �?       @               @      �?      @      �?              �?      @              @                      �?      @     �A@      @      "@      @              @      "@       @      �?      �?              �?      �?              �?      �?              �?       @              @      �?      @               @      �?      �?      �?                      �?              :@      "@     �G@      @       @              �?      @      �?      @              �?      �?              �?      �?              @     �F@       @     �F@       @      2@              1@       @      �?       @                      �?              ;@      �?             �q@     @R@      $@     �B@      $@      "@       @       @      �?      �?      �?                      �?      @      �?              �?      @               @      @       @      @      �?      @      �?                      @      �?                      @              <@     q@      B@     @o@      2@     @o@      1@     @i@      @      :@       @      @       @               @      @              5@              f@      �?     �@@      �?      :@              @      �?      �?      �?      �?                      �?      @             �a@              H@      ,@      H@      *@      :@      $@      8@      @      *@      @      �?      @      �?       @      �?                       @              �?      (@       @      $@               @       @       @      �?              �?       @                      �?      &@               @      @       @                      @      6@      @      @              .@      @              �?      .@       @      .@      �?      @      �?      @                      �?       @                      �?              �?              �?      7@      2@      @      2@      @      ,@      @      @      @               @      @       @                      @              @      �?      @              @      �?      �?              �?      �?              1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��*hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�5         �                    �?�$�����?A           ��@                          �]@"�ZH#��?g           x�@                           �?>a�����?>            �Y@              
             �?#z�i��?            �D@                          �c@д>��C�?             =@                           `@؇���X�?             <@                          @L@������?	             .@                           �?�	j*D�?             *@	       
                   �^@�����H�?             "@������������������������       �                     @              
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @                          �Z@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     �?                           �M@      �?             (@              	            �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @                           �?�]0��<�?&            �N@������������������������       �                    �F@              	             @      �?
             0@������������������������       �        	             ,@������������������������       �                      @       e       	          pff�?�Ç	�X�?)           �|@       <       
             �?�S����?�            `u@        +       	          ����?P��E��?(             R@!       *                    �?�T|n�q�?            �E@"       %                    �?������?             ;@#       $                    e@r�q��?             @������������������������       �                     @������������������������       �                     �?&       )                    h@�����?             5@'       (                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        
             .@������������������������       �                     0@,       ;                    �?>���Rp�?             =@-       4                   �c@      �?             <@.       3                   pm@�KM�]�?	             3@/       2                    @���Q��?             @0       1                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     ,@5       6                    �?X�<ݚ�?             "@������������������������       �                      @7       8                    @K@����X�?             @������������������������       �                     @9       :                    d@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?=       \                   �b@�j�j�?�            �p@>       U       	          ����?P
��M�?�            `n@?       H                    �? 5x ��?�            �j@@       E                    �L@�L���?            �B@A       D                    \@XB���?             =@B       C                   �e@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     7@F       G                    @M@      �?              @������������������������       �                      @������������������������       �                     @I       T                    �O@P����?r             f@J       K                    �?�|���?q             f@������������������������       �        &            �M@L       O                   @[@�T�~~4�?K            @]@M       N                   �l@r�q��?             @������������������������       �                     @������������������������       �                     �?P       Q                   d@ �O�H�?G            �[@������������������������       �        .            �Q@R       S                    �L@�(\����?             D@������������������������       �                    �C@������������������������       �                     �?������������������������       �                     �?V       W                   �Y@ 	��p�?             =@������������������������       �                     �?X       [                   �_@h�����?             <@Y       Z                   �^@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     4@]       b                    �K@�����H�?             ;@^       _                    �? �q�q�?             8@������������������������       �                      @`       a                   0c@      �?	             0@������������������������       �                     �?������������������������       �                     .@c       d       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?f       i                    @D@��|��L�?P            �\@g       h                   �e@؇���X�?             @������������������������       �                     @������������������������       �                     �?j       �                   �r@���B��?L             [@k       v                    �? 9�����?<             V@l       q                   @]@R�}e�.�?             :@m       n                   �^@z�G�z�?             @������������������������       �                     @o       p                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?r       s       
             �?؇���X�?             5@������������������������       �                     .@t       u       	            �?      �?             @������������������������       �                     @������������������������       �                     @w       x       
             �?f���M�?)             O@������������������������       �                     @y       z                    @F@��>4և�?%             L@������������������������       �                     @{       �       
             �?� �	��?!             I@|       }                    �I@*;L]n�?             >@������������������������       �                     @~       �                    @L@�q�����?             9@       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     @�       �                   Pn@ҳ�wY;�?             1@�       �                    �?�eP*L��?             &@������������������������       �                     @�       �                   �b@      �?              @�       �                    @N@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          ����?      �?             4@�       �                     O@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    a@$�q-�?	             *@�       �                     L@�q�q�?             @������������������������       �                     �?�       �                   @d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                   �\@ףp=
�?             4@������������������������       �                     �?�       �                     Q@�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?�       �                    �?<fV���?�            pv@�       �       	          ����?�\��N��?             C@�       �                    �?J�8���?             =@�       �                    �?8�A�0��?             6@������������������������       �                     @�       �                   �_@�\��N��?             3@�       �                   �`@r�q��?             @������������������������       �                     @�       �                   @]@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�n_Y�K�?             *@�       �       	          033�?�q�q�?             (@�       �       	             �?�<ݚ�?             "@�       �                    b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     @�       �                   @`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �       	          ����?�"�����?�            t@�       �                   �i@����!�?.            �T@�       �       
             �?����?�?            �F@������������������������       �                     B@�       �                   0a@�����H�?             "@������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                     P@؀�:M�?            �B@�       �                   �a@      �?             <@�       �                   �^@��Q��?             4@�       �                   �n@؇���X�?             @�       �                    �E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �`@$�q-�?             *@�       �                    �K@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �       	          ����?      �?              @�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                    @xF�8���?�            �m@�       �                   @^@�kb97�?�            �l@�       �                   0m@z�G�z�?            �F@�       �       	             @¦	^_�?             ?@�       �                   @k@$��m��?             :@�       �                    �?���N8�?             5@�       �                    �?�n_Y�K�?             *@�       �       	             �?      �?             $@�       �       
             �?����X�?             @������������������������       �                     �?�       �                   `h@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        
             ,@�       �                    _@0�z��?�?r            @g@�       �                   �[@�C��2(�?             &@������������������������       �                     @�       �                   �\@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                     E@���ib#�?k            �e@������������������������       �                     �?�       �                    �R@�B:�g�?j            �e@������������������������       �        i            �e@������������������������       �                     �?�       �                   �]@      �?              @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       `z@      @      w@     �g@      0@     �U@      ,@      ;@      @      8@      @      8@      @      &@      @      "@      �?       @              @      �?      @      �?                      @      @      �?      @                      �?               @              *@      �?              "@      @      @      @      @                      @      @               @     �M@             �F@       @      ,@              ,@       @              v@     �Y@      r@      K@      =@     �E@      @      B@      @      4@      @      �?      @                      �?       @      3@       @      @              @       @                      .@              0@      6@      @      5@      @      1@       @      @       @      �?       @      �?                       @       @              ,@              @      @       @               @      @              @       @       @               @       @              �?             0p@      &@     `m@       @      j@      @      A@      @      <@      �?      @      �?      @                      �?      7@              @       @               @      @             �e@      @     �e@       @     �M@             �\@       @      @      �?      @                      �?     �[@      �?     �Q@             �C@      �?     �C@                      �?              �?      ;@       @              �?      ;@      �?      @      �?      @                      �?      4@              8@      @      7@      �?       @              .@      �?              �?      .@              �?       @               @      �?             �P@     �H@      �?      @              @      �?             @P@     �E@     �G@     �D@      @      3@      @      �?      @              �?      �?              �?      �?              @      2@              .@      @      @              @      @              D@      6@      @              A@      6@      @              <@      6@      *@      1@              @      *@      (@      @      �?              �?      @              @      &@      @      @      @              @      @      @      �?              �?      @                      @              @      .@      @      @      @              @      @              (@      �?       @      �?      �?              �?      �?      �?                      �?      $@              2@       @              �?      2@      �?      2@                      �?      J@     0s@      4@      2@      3@      $@      *@      "@      @              $@      "@      @      �?      @              �?      �?              �?      �?              @       @      @      @       @      @       @      �?              �?       @                      @      @                      �?      @      �?      @              �?      �?      �?                      �?      �?       @               @      �?              @@     r@      .@     �P@      �?      F@              B@      �?       @               @      �?      @              @      �?              ,@      7@      ,@      ,@      *@      @      �?      @      �?      �?      �?                      �?              @      (@      �?      @      �?              �?      @               @              �?      @      �?      @              @      �?                      �?              "@      1@     �k@      (@     `k@      "@      B@      "@      6@      "@      1@      @      0@      @       @      @      @       @      @              �?       @      @              @       @              @                      @               @      @      �?              �?      @                      @              ,@      @     �f@      �?      $@              @      �?      @      �?                      @       @     �e@      �?              �?     �e@             �e@      �?              @      @              @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ՘�8hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �       
             �?Ly�'^��?B           ��@                           f@�nN@��?B           �@       
       
             �?8$�s���?_            `d@                           �K@     ��?             0@                           �?      �?             @������������������������       �                      @������������������������       �                      @       	                    �?�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@                           �?@9G��?S            `b@              	          ���@@4և���?"             L@                          `X@�X�<ݺ?              K@                           �L@�z�G��?             $@                           �K@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     F@                          c@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?p�C��?1            �V@������������������������       �        &            �R@                           �?�t����?             1@������������������������       �                     (@                           �?���Q��?             @                          �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?        S                   �a@���w��?�            Pu@!       8                    @L@4�d����?�             j@"       7                    �?�q-�?C             Z@#       4       	          ����?㺦���?;            @W@$       3                   �p@�n`���?             ?@%       &                    �E@�z�G��?             4@������������������������       �                      @'       (                    �?�<ݚ�?             2@������������������������       �                     @)       2                    @K@������?
             .@*       +       	             �?8�Z$���?	             *@������������������������       �                     @,       -                   �[@      �?              @������������������������       �                      @.       1                   �m@�q�q�?             @/       0                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@5       6                   �f@0�z��?�?)             O@������������������������       �                     �?������������������������       �        (            �N@������������������������       �                     &@9       R       	          ��� @z�G�z�?I            @Z@:       ?                    �?��C"�b�?:            �T@;       <       	          pff�?����X�?	             ,@������������������������       �                     @=       >                   �\@և���X�?             @������������������������       �                     @������������������������       �                     @@       K                   Ps@�� =[�?1             Q@A       B                   `_@\#r��?,            �N@������������������������       �                      D@C       J                   0a@����X�?             5@D       G                   P`@���Q��?             $@E       F                    �?���Q��?             @������������������������       �                      @������������������������       �                     @H       I       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@L       M                    �O@����X�?             @������������������������       �                     @N       Q       
             �?      �?             @O       P                    �R@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     7@T       y                   �n@�q�q�?W            �`@U       b                    �?j���� �?,             Q@V       ]                    c@���Q��?             9@W       X                    �?�	j*D�?             *@������������������������       �                      @Y       Z       	          ����?z�G�z�?             @������������������������       �                      @[       \       	          hff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @^       _                   �l@�8��8��?             (@������������������������       �                     $@`       a                   �m@      �?              @������������������������       �                     �?������������������������       �                     �?c       n                   ``@�^�����?            �E@d       g       
             �?�8��8��?             8@e       f       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?h       i       	          ����?P���Q�?             4@������������������������       �                     "@j       m                   �b@�C��2(�?	             &@k       l                   �m@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @o       p       
             �?D�n�3�?             3@������������������������       �                     @q       t                    �?     ��?	             0@r       s                   �b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?u       x       	          pff�?�C��2(�?             &@v       w                   `c@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @z       �                   u@     ��?+             P@{       |                    �I@�X�C�?&             L@������������������������       �                     4@}       �                    �?      �?             B@~                          p@�z�G��?             >@������������������������       �                     "@�       �       	          `ff�?և���X�?             5@�       �                   pc@���Q��?
             .@�       �                    �?���!pc�?             &@�       �       	             �?�����H�?             "@������������������������       �                     @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @������������������������       �                      @�       �                    �L@�@��T�?            �y@�       �                    I@��[��^�?�            0t@�       �       	            �?��2(&�?             6@�       �                    @I@���Q��?             @�       �                   @b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        
             1@�       �                    �?t���W�?�            �r@�       �                   �a@�<ݚ�?+             R@�       �       	          433�?h�����?             <@������������������������       �                     8@�       �                   �r@      �?             @������������������������       �                      @�       �                   `b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�X���?             F@������������������������       �                     $@�       �                    �D@�ʻ����?             A@������������������������       �                      @�       �                    o@R�}e�.�?             :@�       �       	          ����?      �?
             0@�       �                    ]@@4և���?             ,@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �`@      �?             $@�       �                   �e@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    @L@0<�q �?�            �l@�       �                    �?0���|�?�             l@�       �                    �J@ףp=
�?             >@�       �                   �]@`2U0*��?             9@�       �                   �d@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@�       �                    �?���Q��?             @�       �                   `f@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                   @n@@�����?r            `h@������������������������       �        M            �`@�       �                    �?��v$���?%            �N@������������������������       �                    �F@�       �                   �b@      �?	             0@������������������������       �                      @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   `Q@��+�ޯ�??            �V@�       �                    �?z�G�z�?             4@�       �                   �^@և���X�?             @������������������������       �                     �?�       �                   `_@�q�q�?             @�       �                    �P@�q�q�?             @�       �                   �V@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        	             *@�       �                    �?��W3�?/            �Q@�       �       	            �?��
P��?            �A@�       �                    ]@��+7��?             7@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �b@r�q��?
             2@�       �                   Pc@��S�ۿ?             .@������������������������       �                     &@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�8��8��?             (@�       �       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                    �M@�<ݚ�?             B@�       �                    @���Q��?             $@�       �       	          833@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   `c@r�q��?             @�       �                    @M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�                         ht@$�q-�?             :@�       �                    �? �q�q�?             8@������������������������       �                     3@�       �                    �?z�G�z�?             @������������������������       �                      @                         @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?�t�b�7     h�h(h+K ��h-��R�(KMKK��h_�BP       �z@     �~@      W@     �y@      "@     @c@      @      *@       @       @       @                       @      �?      &@      �?                      &@      @     �a@      @      J@      @     �I@      @      @      @      @              @      @                      @              F@      �?      �?              �?      �?               @     @V@             �R@       @      .@              (@       @      @       @       @               @       @                      �?     �T@      p@      <@     �f@      @     @X@      @     �U@      @      9@      @      ,@       @              @      ,@              @      @      &@       @      &@              @       @      @               @       @      @      �?      @      �?                      @      �?               @                      &@      �?     �N@      �?                     �N@              &@      5@      U@      5@     �N@      $@      @      @              @      @              @      @              &@     �L@      @     �K@              D@      @      .@      @      @       @      @       @                      @      @      �?      @                      �?              &@      @       @      @               @       @       @      �?              �?       @                      �?              7@     �K@     @S@      D@      <@      $@      .@      "@      @       @              �?      @               @      �?       @      �?                       @      �?      &@              $@      �?      �?      �?                      �?      >@      *@      6@       @      @      �?      @                      �?      3@      �?      "@              $@      �?      @      �?      @                      �?      @               @      &@      @              @      &@      @      �?      @                      �?      �?      $@      �?      @              @      �?                      @      .@     �H@      "@     �G@              4@      "@      ;@      "@      5@              "@      "@      (@      "@      @       @      @       @      �?      @               @      �?              �?       @                       @      �?      @      �?                      @              @              @      @       @      @                       @     �t@     �T@     �q@     �D@      @      3@      @       @      �?       @      �?                       @       @                      1@     pq@      6@      L@      0@      ;@      �?      8@              @      �?       @              �?      �?              �?      �?              =@      .@      $@              3@      .@               @      3@      @      ,@       @      *@      �?      �?      �?              �?      �?              (@              �?      �?              �?      �?              @      @       @      @              @       @              @             �k@      @     �k@      @      ;@      @      8@      �?      @      �?              �?      @              4@              @       @       @       @       @                       @      �?             @h@      �?     �`@              N@      �?     �F@              .@      �?       @              @      �?              �?      @               @       @      �?       @               @      �?              �?              I@     �D@      @      0@      @      @              �?      @       @      �?       @      �?      �?              �?      �?                      �?      @                      *@      G@      9@      2@      1@      1@      @       @      @              @       @              .@      @      ,@      �?      &@              @      �?              �?      @              �?       @      �?                       @      �?      &@      �?      �?              �?      �?                      $@      <@       @      @      @      @      �?      @                      �?      �?      @      �?       @      �?                       @              @      8@       @      7@      �?      3@              @      �?       @               @      �?              �?       @              �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�4hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKh~�BH4         �                    �?�7i���?I           ��@       E                    �?j�	k�?X           �@       6       	          ����?�萻/#�?~             i@              
             �?��/���?b             d@              	          833�?����?/            �S@������������������������       �                     G@                          �r@     ��?             @@                          �[@8�A�0��?             6@	                          p@����X�?             @
                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @                           �?������?             .@                          �_@���|���?             &@������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@                          `X@rp��P��?3            �T@������������������������       �                     @       3                    �?�G�z.�?2             T@       0                    �?     ��?(             P@                           �?�1�`jg�?#            �K@������������������������       �                     @       #                    �?`�Q��?             I@                            G@���|���?             &@������������������������       �                     @                            �L@�q�q�?             @������������������������       �                     @!       "                   p`@�q�q�?             @������������������������       �                      @������������������������       �                     �?$       +                    b@�θ�?            �C@%       &                    �I@      �?             @@������������������������       �                     4@'       *                    c@�q�q�?	             (@(       )                   @E@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     @,       -                   `Y@����X�?             @������������������������       �                     �?.       /                   �s@r�q��?             @������������������������       �                     @������������������������       �                     �?1       2                   @[@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @4       5                    U@      �?
             0@������������������������       �                     �?������������������������       �        	             .@7       B                    �Q@ףp=
�?             D@8       ?                    �?�˹�m��?             C@9       <                   pd@z�G�z�?             $@:       ;                   Pe@      �?              @������������������������       �                     �?������������������������       �                     �?=       >                    �O@      �?              @������������������������       �                     @������������������������       �                     �?@       A                   Pd@h�����?             <@������������������������       �                     ;@������������������������       �                     �?C       D       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?F       I                    Z@�X�R�?�            @u@G       H       
             �?�����?             3@������������������������       �        	             *@������������������������       �                     @J       o       
             �?�����?�            t@K       h       	          ���@8�A�0��?9             V@L       O                   �[@      �?3             T@M       N                    �?      �?              @������������������������       �                     �?������������������������       �                     @P       Y                    �?�E����?-             R@Q       R                    a@\-��p�?             =@������������������������       �                     .@S       X                   �c@����X�?             ,@T       U                    �P@�C��2(�?             &@������������������������       �                      @V       W                   @`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @Z       a       	          ����?�+��<��?            �E@[       `                   @_@�����?             3@\       _                   �e@      �?              @]       ^                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@b       g                   �c@      �?             8@c       d                    �?"pc�
�?             6@������������������������       �                     "@e       f       	          `ff�?�	j*D�?	             *@������������������������       �                     "@������������������������       �                     @������������������������       �                      @i       n       	          ���@      �?              @j       k                    �?؇���X�?             @������������������������       �                     @l       m                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?p       �                    �Q@�t M\�?�             m@q       �                   h@p�|�i�?�            �l@r       {                    �?���{h�?�            `l@s       t                    @L@ qP��B�?T             `@������������������������       �        I             ]@u       v                   �_@�θ�?             *@������������������������       �                     �?w       z                    �?r�q��?
             (@x       y                   pb@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@|       �                   pf@ؗp�'ʸ?=            �X@}       �                   �`@`�q�0ܴ?9            �W@~       �                    �L@�:�]��?            �I@       �                    d@���7�?             F@�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   0n@�(\����?             D@������������������������       �                     9@�       �                   �n@��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@�       �                    @����X�?             @�       �                   �d@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �E@�       �                   �`@      �?             @�       �                    �F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       
             �?�&�ѩ��?�            �w@�       �                    �R@     ��?�             t@�       �                   Pe@���.n�?�            �s@�       �                   pa@(�5�f��?5            �S@������������������������       �        3             S@������������������������       �                     @�       �                    �?x��)f��?�            `m@�       �                   pb@ �M*k�?}            �h@�       �                    f@ ,��-�?q             f@�       �                   �e@�}�+r��?n            `e@������������������������       �                     �?�       �                   j@Pq�����?m            @e@�       �                   �i@"pc�
�?             6@�       �       	          ����?�����H�?             2@������������������������       �                     "@�       �                   `i@�<ݚ�?             "@�       �       
             �?�q�q�?             @������������������������       �                     @�       �                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   @\@      �?             @������������������������       �                      @������������������������       �                      @�       �       	          ����?�?�|�?\            �b@�       �                    �?      �?	             (@������������������������       �                      @�       �                     P@�z�G��?             $@�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   �[@�|�l�?S             a@�       �                   �m@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �        K             _@�       �                   `^@      �?             @������������������������       �                      @�       �       	          433@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �a@z�G�z�?             4@�       �                    �?���Q��?             $@������������������������       �                      @�       �       	          `ff�?      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@�       �                    �?P����?             C@�       �                   Pm@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��a�n`�?             ?@�       �       	             �?�X����?             6@�       �                    �?���|���?             &@������������������������       �                     @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                     "@�       �       	             @      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?�\��N��?'            �L@�       �                    �?      �?             D@������������������������       �                     @�       �                   ``@��G���?            �B@�       �                    �?�IєX�?             1@������������������������       �                     &@�       �                    _@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?�z�G��?             4@�       �                    h@      �?              @�       �                   @b@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @M@�8��8��?             (@������������������������       �                     $@�       �                    @N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     1@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       pz@     �~@     �v@     �f@      U@     @]@      T@     @T@      3@     �M@              G@      3@      *@      "@      *@      @       @      �?       @      �?                       @      @              @      &@      @      @              @      @       @               @      @                      @      $@             �N@      6@              @     �N@      3@      G@      2@     �C@      0@      @              A@      0@      @      @              @      @       @      @              �?       @               @      �?              >@      "@      <@      @      4@               @      @       @      �?              �?       @                      @       @      @      �?              �?      @              @      �?              @       @               @      @              .@      �?              �?      .@              @      B@      @     �A@       @       @      �?      �?              �?      �?              �?      @              @      �?              �?      ;@              ;@      �?              �?      �?              �?      �?             Pq@     �O@      @      *@              *@      @             �p@      I@      J@      B@      I@      >@      �?      @      �?                      @     �H@      7@      9@      @      .@              $@      @      $@      �?       @               @      �?       @                      �?              @      8@      3@      @      *@      @       @      @      �?      @                      �?              �?              &@      2@      @      2@      @      "@              "@      @      "@                      @               @       @      @      �?      @              @      �?       @      �?                       @      �?             `k@      ,@     `k@      "@     `k@       @     �_@      @      ]@              $@      @              �?      $@       @      �?       @      �?                       @      "@             @W@      @     �V@      @     �G@      @      E@       @      @      �?              �?      @             �C@      �?      9@              ,@      �?              �?      ,@              @       @      @      �?      @                      �?              �?     �E@              @      �?      �?      �?      �?                      �?       @                      �?              @      O@     �s@     �A@     �q@      @@     �q@      @      S@              S@      @              =@     �i@      0@     �f@      (@     �d@      "@     @d@      �?               @     @d@      @      2@       @      0@              "@       @      @       @      @              @       @      �?              �?       @                      @       @       @       @                       @      @      b@      @      "@               @      @      @      @      @              @      @                      @      �?     �`@      �?      &@      �?                      &@              _@      @      @               @      @      �?      @                      �?      @      0@      @      @       @               @      @              @       @      �?       @                      �?              $@      *@      9@      @      �?      @                      �?      @      8@      @      .@      @      @              @      @      �?              �?      @                      &@              "@      @      @      @                      @      ;@      >@      $@      >@      @              @      >@      �?      0@              &@      �?      @              @      �?              @      ,@      @      @      �?      @               @      �?      �?              �?      �?              @              �?      &@              $@      �?      �?      �?                      �?      1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�BX7         �       
             �?TU�`��?@           ��@       Y                    �?2�!	s��?U           Ѐ@       V                   �e@7~���?�            x@                           �?�x+M���?�            �w@                          �_@�{��?��?"             K@                          �r@      �?             0@                            G@�θ�?	             *@������������������������       �                     �?	       
                   @_@r�q��?             (@������������������������       �                      @������������������������       �                     $@������������������������       �                     @                           �?�?�'�@�?             C@              
             �?      �?
             0@������������������������       �                     @                           �?r�q��?             (@                           b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @              	          033�?��2(&�?             6@������������������������       �                     $@                           `@      �?             (@������������������������       �                     @              	          033�?և���X�?             @������������������������       �                     @������������������������       �                     @                          �U@��8=��?�            �t@������������������������       �                      @       C                   pb@�@�?�            `t@       "                   �Q@�B𛇯?�            �q@        !       	          033�?      �?             @������������������������       �                     @������������������������       �                     �?#       $       	          433�?`�X$��?�            pq@������������������������       �        %             M@%       :                   ``@X�t3�ܱ?�            �k@&       1                    �?��Wv��?C             [@'       (       	             �?�J�4�?             9@������������������������       �                     �?)       0       	             �?      �?             8@*       /                    �?d}h���?	             ,@+       .       	          033�?�q�q�?             "@,       -                   8q@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@2       9                    �L@P��BNֱ?5            �T@3       8                    \@0G���ջ?              J@4       7                   pp@z�G�z�?
             .@5       6                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     $@������������������������       �                    �B@������������������������       �                     ?@;       B                    �K@�H�I���?F            @\@<       =                    @K@`���i��?             F@������������������������       �                     B@>       A                   �n@      �?              @?       @                   �k@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        +            @Q@D       I                   �b@�T|n�q�?            �E@E       F       	          433�?�q�q�?             @������������������������       �                      @G       H                   l@      �?             @������������������������       �                      @������������������������       �                      @J       K                   �b@�L���?            �B@������������������������       �                     0@L       S                   �r@؇���X�?             5@M       N                     L@�KM�]�?             3@������������������������       �        	             *@O       P                    �?�q�q�?             @������������������������       �                      @Q       R                    �?      �?             @������������������������       �                      @������������������������       �                      @T       U                    x@      �?              @������������������������       �                     �?������������������������       �                     �?W       X       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @Z       m                   �h@��7�G%�?e             c@[       ^                    @J@t/*�?            �G@\       ]                    �?�}�+r��?             3@������������������������       �                     �?������������������������       �        
             2@_       l                   �e@      �?             <@`       k                   �c@�J�4�?             9@a       j       	          033�?      �?             8@b       c       
             �?d}h���?	             ,@������������������������       �                      @d       i                    Z@�8��8��?             (@e       f                    �?      �?             @������������������������       �                      @g       h                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     �?������������������������       �                     @n                          �a@~|z����?G            �Z@o       v                   pm@@�0�!��?             A@p       q                    @K@�q�q�?
             (@������������������������       �                      @r       u                   @l@z�G�z�?             $@s       t                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?w       x                   �r@�C��2(�?             6@������������������������       �        	             .@y       ~                    @����X�?             @z       }                   �t@r�q��?             @{       |                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    @L@<ݚ)�?/             R@�       �                   Xp@ s�n_Y�?!             J@�       �                    �?�KM�]�?             C@�       �                   �`@�L���?            �B@�       �                    �?�IєX�?             A@�       �                   �d@XB���?             =@������������������������       �                     0@�       �       
             �?$�q-�?             *@�       �                   �\@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @J@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   Hr@      �?
             ,@�       �                    �?�<ݚ�?             "@�       �                    �?���Q��?             @�       �                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       	          `ff @�G�z��?             4@�       �                   �l@����X�?             ,@������������������������       �                      @�       �       	          ����?r�q��?	             (@�       �                   `d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    o@ףp=
�?             $@�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   pa@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�[%�r�?�            �w@�       �                   �]@r�q��?M             ^@�       �                    �J@�q�q�?             >@�       �                   �a@��.k���?
             1@������������������������       �                     @�       �                    @F@���!pc�?             &@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �P@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?�       �                   �c@b�2�tk�?;            �V@�       �       	          `ff�?l��
I��?             ;@�       �                   �_@�+e�X�?             9@�       �       	             �?$�q-�?             *@�       �                   �]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�       �                   �b@�q�q�?             (@�       �                    �?�<ݚ�?             "@�       �                   @E@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?�w��@�?+            �O@�       �                   d@���7�?             F@������������������������       �                    �A@�       �                   �q@�<ݚ�?             "@�       �                   @d@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   `_@�d�����?             3@������������������������       �                      @�       �                    �?@�0�!��?             1@������������������������       �                     &@�       �                    @I@      �?             @������������������������       �                     @������������������������       �                     @�       �                   0h@����?�            @p@�       �                   �_@ T[����?�            p@�       �                   �c@"pc�
�?            �@@������������������������       �                     @�       �                    �? 	��p�?             =@�       �                    @ 7���B�?             ;@������������������������       �                     8@�       �                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �P@      �?�             l@�       �                   0`@���!pc�?             &@�       �                    @H@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    @M@���~qޢ?�            �j@�       �                   @[@�eGk�T�?r            �g@�       �                    �?r�q��?	             (@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                      @�       �                   `m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        i            @f@�       �                   ps@���}<S�?             7@�       �                    �M@P���Q�?             4@�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             0@�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       @y@     �@     �W@     �{@      ?@      v@      =@     v@      &@     �E@      @      $@      @      $@      �?               @      $@       @                      $@      @              @     �@@       @      ,@              @       @      $@       @       @       @                       @               @      @      3@              $@      @      "@              @      @      @      @                      @      2@     `s@       @              0@     `s@      "@      q@      �?      @              @      �?               @     �p@              M@       @     �j@      @     @Y@      @      5@      �?              @      5@      @      &@      @      @       @      @              @       @              �?                      @              $@      @      T@      @     �H@      @      (@      @       @               @      @                      $@             �B@              ?@      �?      \@      �?     �E@              B@      �?      @      �?      @              @      �?                      @             @Q@      @      B@      @       @       @               @       @       @                       @      @      A@              0@      @      2@       @      1@              *@       @      @               @       @       @       @                       @      �?      �?      �?                      �?       @      �?              �?       @              P@     @V@       @     �C@      �?      2@      �?                      2@      @      5@      @      5@      @      5@      @      &@       @              �?      &@      �?      @               @      �?      �?      �?                      �?               @              $@      �?              @              L@      I@      @      <@      @       @       @               @       @      �?       @      �?                       @      �?               @      4@              .@       @      @      �?      @      �?      �?      �?                      �?              @      �?              I@      6@     �D@      &@      A@      @      A@      @      @@       @      <@      �?      0@              (@      �?      @      �?              �?      @              @              @      �?      @                      �?       @      �?       @                      �?              �?      @      @       @      @       @      @       @      �?       @                      �?               @              @      @              "@      &@      @      $@       @               @      $@      �?      �?      �?                      �?      �?      "@      �?       @               @      �?                      @      @      �?              �?      @             Ps@     �Q@     @P@     �K@      $@      4@      "@       @      @              @       @              @      @       @      @                       @      �?      (@              (@      �?             �K@     �A@       @      3@      @      3@      �?      (@      �?      �?      �?                      �?              &@      @      @       @      @       @      @              @       @                      @      @               @             �G@      0@      E@       @     �A@              @       @      @      �?              �?      @                      �?      @      ,@       @              @      ,@              &@      @      @      @                      @     �n@      0@     �n@      *@      ;@      @              @      ;@       @      :@      �?      8@               @      �?       @                      �?      �?      �?              �?      �?              k@      @       @      @      @      @      @                      @      @              j@      @     �g@       @      $@       @      @              @       @       @              �?       @      �?                       @     @f@              5@       @      3@      �?      @      �?      @                      �?      0@               @      �?              �?       @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��1zhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK녔h~�Bh3         �                    �?\r��ۖ�?A           ��@       A                    �?�!��CG�?4           �@                          0a@ڡR����?            �h@                           �?�U�=���?*            �P@       
                    �?X�Cc�?             ,@              
             �?���|���?             &@������������������������       �                     @       	                   �^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @              
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     J@       &       
             �?
j*D>�?U            @`@              	             �?     ��?'             P@              	          833�?~�4_�g�?             F@������������������������       �                     .@                          `]@J�8���?             =@������������������������       �                     @                          Pr@�q�q�?             8@              	          ����?     ��?
             0@                           @I@�����H�?             "@                           b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @        %                    _@P���Q�?             4@!       "                   �r@�����H�?             "@������������������������       �                     @#       $                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@'       (                   �b@r�q��?.            �P@������������������������       �                     A@)       *                   @c@     ��?             @@������������������������       �                      @+       <                    b@�z�G��?             >@,       5                   �_@z�G�z�?             9@-       .                   �c@      �?              @������������������������       �                      @/       4                   0k@�q�q�?             @0       1                    �?      �?             @������������������������       �                     �?2       3                     I@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @6       ;                    �?�IєX�?             1@7       :                    �?z�G�z�?             @8       9                    �M@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@=       @                    �I@z�G�z�?             @>       ?                   `m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @B       }                    �?�Rez��?�            �s@C       x                   Pd@��g�g�?�            �m@D       o       
             �?$�b���?�            `l@E       `       	          ����?�][�M_�?u            `h@F       G                   �i@H�V�e��?&             Q@������������������������       �                     @@H       [                   �a@b�2�tk�?             B@I       J                    �?
;&����?             7@������������������������       �                     �?K       N                    �?�eP*L��?             6@L       M                    �D@      �?             @������������������������       �                      @������������������������       �                      @O       V                    n@X�<ݚ�?
             2@P       U                     P@"pc�
�?             &@Q       T                     J@ףp=
�?             $@R       S                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?W       Z       	          433�?؇���X�?             @X       Y       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @\       _                   @e@8�Z$���?             *@]       ^                   �n@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?a       h                   �a@�U���?O            �_@b       g       	          ����?���1��?C            �Z@c       d                   @_@ 7���B�?             ;@������������������������       �                     7@e       f                   �i@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        0             T@i       l       
             �?ףp=
�?             4@j       k                    U@      �?             @������������������������       �                     �?������������������������       �                     @m       n                   �Z@      �?	             0@������������������������       �                     �?������������������������       �                     .@p       w                   �`@      �?             @@q       v                   �r@��.k���?             1@r       s                   �[@��S���?	             .@������������������������       �                     @t       u                     P@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@y       |                   xs@X�<ݚ�?             "@z       {       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @~                          0a@�}�+r��?)             S@������������������������       �                    �B@�       �       	          `ff�?��-�=��?            �C@�       �                   `c@      �?             @������������������������       �                     @������������������������       �                     @�       �                   @s@Pa�	�?            �@@������������������������       �                     ?@�       �                   `t@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �`@~j�$s�?           �y@�       �       
             �?��
ц��?S            @`@�       �                   @^@>A�F<�?/             S@�       �                    �? �o_��?             I@�       �                    �?����X�?             @�       �                   `X@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    @L@RB)��.�?            �E@�       �                    �?��
ц��?             *@�       �       	             �?�z�G��?             $@�       �                   `X@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	             �?ףp=
�?             >@������������������������       �                     2@�       �                    �?      �?             (@������������������������       �                     @������������������������       �                     "@������������������������       �                     :@�       �                    �P@PN��T'�?$             K@�       �                   �c@=QcG��?             �G@�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                    �D@�       �                    �?����X�?             @������������������������       �                     �?�       �                    @r�q��?             @�       �                     R@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    I@h�d.��?�            �q@�       �                   �a@�q�q�?             "@������������������������       �                      @�       �                    @؇���X�?             @�       �                    �?z�G�z�?             @������������������������       �                     @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @L@֙S}o�?�            �p@�       �                   �l@l}N+V5�?�            �h@�       �       
             �?���N8�?D            @Z@�       �                    �?X�Cc�?             ,@�       �                   �c@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �e@      �?              @������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        8            �V@�       �       
             �?Ʋ(>^�?@            @W@�       �                   0a@`՟�G��?             ?@�       �                    ]@`�Q��?             9@������������������������       �                     @�       �                    @R���Q�?             4@�       �                   hp@�KM�]�?             3@������������������������       �                     ,@�       �                    �?���Q��?             @������������������������       �                      @�       �                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        .             O@�       �                    �?���o,��?.            @R@�       �       
             �?��.k���?             A@�       �                   �o@�E��ӭ�?             2@������������������������       �                     @�       �                    q@�eP*L��?             &@������������������������       �                     @�       �                    `P@      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �M@     ��?	             0@�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@�       �                    @O@8�Z$���?            �C@�       �                   �`@�+e�X�?             9@�       �       	          @33�?�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �        
             0@������������������������       �        	             ,@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       py@     �@     �\@     �x@      T@      ]@      @     �N@      @      "@      @      @              @      @      �?              �?      @              �?       @      �?                       @              J@     �R@     �K@      4@      F@      3@      9@              .@      3@      $@              @      3@      @      &@      @       @      �?       @      �?       @                      �?      @              @      @      @                      @       @              �?      3@      �?       @              @      �?      �?      �?                      �?              &@     �K@      &@      A@              5@      &@               @      5@      "@      4@      @      @      @               @      @       @       @       @              �?       @      �?       @                      �?       @              0@      �?      @      �?      @      �?      @                      �?      �?              (@              �?      @      �?      �?              �?      �?                      @      A@     `q@      >@     �i@      9@     @i@      1@     @f@      ,@      K@              @@      ,@      6@      (@      &@              �?      (@      $@       @       @               @       @              $@       @      "@       @      "@      �?       @      �?              �?       @              @                      �?      �?      @      �?      �?              �?      �?                      @       @      &@      �?      &@      �?                      &@      �?              @      _@      �?     �Z@      �?      :@              7@      �?      @      �?                      @              T@       @      2@      �?      @      �?                      @      �?      .@      �?                      .@       @      8@       @      "@       @      @              @       @      �?       @                      �?               @              .@      @      @       @      @       @                      @      @              @      R@             �B@      @     �A@      @      @      @                      @      �?      @@              ?@      �?      �?      �?                      �?     Pr@     @]@      N@     �Q@      ,@      O@      ,@      B@      @       @      @      �?              �?      @                      �?      "@      A@      @      @      @      @      @      @      @                      @              @      @              @      ;@              2@      @      "@      @                      "@              :@      G@       @      F@      @      @      @      @                      @     �D@               @      @      �?              �?      @      �?       @      �?                       @              @      m@     �G@      @      @       @              �?      @      �?      @              @      �?      �?      �?                      �?               @     �l@     �D@     `f@      3@      Y@      @      "@      @      @      �?              �?      @              @      @               @      @       @      @              �?       @      �?                       @     �V@             �S@      ,@      1@      ,@      1@       @              @      1@      @      1@       @      ,@              @       @       @              �?       @      �?                       @              �?              @      O@             �I@      6@      2@      0@      @      *@              @      @      @      @               @      @              @       @      �?       @                      �?      *@      @      �?      @              @      �?              (@             �@@      @      3@      @      @      @      @                      @      0@              ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJT�bhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�;         �                    �?�ܢ����?N           ��@       �                    �?��-�7k�?a           `�@       r       	          033�?tk~X���?            {@                           �?<�hgێ�?�            �x@              
             �?�X�<ݺ?P            �_@                           @C@     ��?             @@������������������������       �                     �?       	                    �G@��� ��?             ?@������������������������       �                     "@
                           b@"pc�
�?             6@                          @q@ףp=
�?             4@������������������������       �        
             *@                           �?����X�?             @������������������������       �                     @                           _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �?`Ql�R�?9            �W@                          d@ףp=
�?             $@������������������������       �                      @                          �q@      �?              @������������������������       �                     �?������������������������       �                     �?                            R@ ��N8�?1             U@������������������������       �        0            �T@������������������������       �                     �?       C       
             �?@�h�|5�?�            �p@       *                    �?v�_���?3            �S@       )                    �?�d�����?             C@       "                     M@      �?             @@        !                   �e@`2U0*��?             9@������������������������       �                     8@������������������������       �                     �?#       $       	          ����?և���X�?             @������������������������       �                      @%       &                    �N@���Q��?             @������������������������       �                      @'       (       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @+       >                   `o@v�2t5�?            �D@,       1                    �?��H�}�?             9@-       0                   `Y@ףp=
�?             $@.       /                   @_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @2       5                    �?��S���?             .@3       4                    @L@      �?              @������������������������       �                     @������������������������       �                     @6       7                    \@����X�?             @������������������������       �                      @8       =                   �`@���Q��?             @9       :                    �L@�q�q�?             @������������������������       �                     �?;       <                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @?       B                   Pq@      �?	             0@@       A       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@D       W                    @L@�*/�8V�?w            �g@E       L                    �? sAr�=�?[            �b@F       I                   i@�t����?             1@G       H                    @A@�q�q�?             @������������������������       �                      @������������������������       �                     @J       K                   `e@�C��2(�?
             &@������������������������       �        	             $@������������������������       �                     �?M       N                    �I@ ����O�?M            ``@������������������������       �        2            @V@O       R                    @J@�����?             E@P       Q                    �?d}h���?             ,@������������������������       �                     @������������������������       �                     &@S       T                    �?h�����?             <@������������������������       �                     4@U       V                   �[@      �?              @������������������������       �                     �?������������������������       �                     @X       q                    �?��Q���?             D@Y       b                    �?">�֕�?            �A@Z       a       	          @33�?z�G�z�?             $@[       `                    @�<ݚ�?             "@\       ]                   0c@      �?              @������������������������       �                     @^       _                   �e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?c       n       	             �?��H�}�?             9@d       m       	          ����?����X�?             5@e       f                   �a@ҳ�wY;�?             1@������������������������       �                     $@g       l                     @؇���X�?             @h       k       	          @33�?      �?             @i       j                   `a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @o       p                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @s       �                    @�q�q�?            �C@t       �                   �`@r٣����?            �@@u       �       
             �?      �?
             0@v       }                    �N@�q�q�?             (@w       |                   `o@؇���X�?             @x       y                   @_@�q�q�?             @������������������������       �                     �?z       {                   pi@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @~                          �\@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             1@�       �                   `U@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    _@f���M�?O             _@�       �                   �c@�&=�w��?"            �J@������������������������       �                    �F@�       �                   0d@      �?              @������������������������       �                      @������������������������       �                     @�       �       
             �?DX�\��?-            �Q@�       �                    �J@z�G�z�?            �A@�       �                   f@�q�q�?             (@�       �                   j@�z�G��?             $@������������������������       �                      @�       �                   `@      �?              @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �x@���}<S�?             7@�       �                    @���7�?             6@������������������������       �                     3@�       �                    @P@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �L@������?             B@������������������������       �                     8@�       �                    @M@�8��8��?	             (@�       �                   �a@�q�q�?             @������������������������       �                     �?�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   �b@������?�            �v@�       �                    @�KM�]�?�            0t@�       �       	          ����?�ʠ����?�            t@�       �                    �N@���-T��?|            @g@�       �       
             �?:��o#@�?_            �a@�       �                   `f@x���� �?R             ^@�       �       	          hff�?�y��*�?O             ]@������������������������       �                     >@�       �                   �n@�T|n�q�?:            �U@�       �                    �?��$�4��?(            �M@������������������������       �                     @�       �                   �\@      �?#             J@�       �                     E@�q�q�?             @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	          033�?�3Ea�$�?             G@�       �                   �i@      �?             @������������������������       �                      @������������������������       �                      @�       �       	          033�?r�q��?             E@�       �                    �?��� ��?             ?@������������������������       �                     �?�       �                    �?ףp=
�?             >@�       �                    @L@�8��8��?             8@������������������������       �        
             0@�       �                   �`@      �?              @�       �                   �Y@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?���!pc�?             &@�       �                    �C@�q�q�?             "@������������������������       �                     @�       �                   �h@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �L@ 7���B�?             ;@������������������������       �                     9@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    w@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?և���X�?             5@�       �       	             �?���Q��?
             .@������������������������       �                     @�       �                   �`@      �?              @�       �                    �?      �?             @�       �                    @M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    \@����?�?            �F@�       �                   @Z@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     D@�       �                    �R@`Ӹ����?X            �`@�       �                   @^@��ɉ�?U            @`@�       �                   @M@r�q��?             8@�       �                    @N@և���X�?             @�       �                    �I@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�IєX�?             1@�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             .@������������������������       �        F            �Z@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�                          �?�q�q�?            �C@                          �?�q�����?             9@                         @D@؇���X�?             @������������������������       �                     �?������������������������       �                     @                         �?�q�q�?             2@������������������������       �                     @                         @K@؇���X�?
             ,@������������������������       �                      @      	                   _@�q�q�?             @������������������������       �                     �?
                        �c@���Q��?             @������������������������       �                     �?            
             �?      �?             @������������������������       �                     �?                        �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@�t�b�h     h�h(h+K ��h-��R�(KMKK��h_�B       �z@     p~@     0w@      g@     pt@     @Z@     �s@     �S@     �]@      @      ;@      @              �?      ;@      @      "@              2@      @      2@       @      *@              @       @      @              �?       @      �?                       @               @      W@       @      "@      �?       @              �?      �?      �?                      �?     �T@      �?     �T@                      �?     `h@      R@      ;@      J@      $@      <@      @      <@      �?      8@              8@      �?              @      @               @      @       @       @              �?       @      �?                       @      @              1@      8@      0@      "@      "@      �?       @      �?              �?       @              @              @       @      @      @      @                      @       @      @               @       @      @       @      �?      �?              �?      �?              �?      �?                       @      �?      .@      �?      @      �?                      @              &@      e@      4@     `a@      "@      (@      @       @      @       @                      @      $@      �?      $@                      �?     �_@      @     @V@              C@      @      &@      @              @      &@              ;@      �?      4@              @      �?              �?      @              =@      &@      8@      &@       @       @      @       @      @      �?      @              �?      �?              �?      �?                      �?      �?              0@      "@      .@      @      &@      @      $@              �?      @      �?      @      �?      �?      �?                      �?               @              @      @              �?      @              @      �?              @              *@      :@       @      9@       @       @      @      @      �?      @      �?       @              �?      �?      �?              �?      �?                      @      @      �?              �?      @              @      �?      @                      �?              1@      @      �?              �?      @              F@      T@       @     �I@             �F@       @      @       @                      @      E@      =@      @      <@      @      @      @      @       @              �?      @      �?      �?              �?      �?                      @       @               @      5@      �?      5@              3@      �?       @               @      �?              �?             �A@      �?      8@              &@      �?       @      �?      �?              �?      �?      �?                      �?      "@              N@     �r@      A@     r@     �@@      r@      ;@     �c@      :@     �\@      1@     �Y@      ,@     �Y@              >@      ,@      R@      *@      G@              @      *@     �C@      @       @              �?      @      �?      @                      �?      "@     �B@       @       @               @       @              @     �A@      @      ;@      �?              @      ;@       @      6@              0@       @      @       @      @              @       @                      @      �?      @              @      �?              @       @      @      @              @      @      @      @                      @               @      �?      :@              9@      �?      �?              �?      �?              @      �?      @                      �?      "@      (@      "@      @      @               @      @       @       @      �?       @               @      �?              �?                      @              @      �?      F@      �?      @              @      �?                      D@      @      `@      @     �_@      @      4@      @      @      @      �?              �?      @                      @      �?      0@      �?      �?      �?                      �?              .@             �Z@       @      @              @       @              �?      �?              �?      �?              :@      *@      (@      *@      @      �?              �?      @              @      (@      @               @      (@               @       @      @              �?       @      @      �?              �?      @              �?      �?       @               @      �?              ,@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��	hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�>         �                    �?�7i���?C           ��@       e                   �`@��I(���?�           H�@                          `[@�t����?�            r@                           �?B�1V���?>            @X@                            J@r�q��?             8@������������������������       �                     @                           �?ҳ�wY;�?             1@       	       
             �?d}h���?
             ,@������������������������       �                     $@
                           �?      �?             @������������������������       �                      @                           @M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           [@��pBI�?-            @R@������������������������       �                     �?                           �O@�k~X��?,             R@������������������������       �        !            �J@              	          433�?�}�+r��?             3@                          �X@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@       &                    �?r�q��?�             h@              	          ����?H�V�e��?             A@                           �P@���}<S�?             7@������������������������       �        
             4@                          �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @        !                    @M@�eP*L��?             &@������������������������       �                     @"       %                    �?؇���X�?             @#       $                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @'       P       
             �?n��s�Z�?p            �c@(       C                    �?�y��*�?Q             ]@)       *       
             �?�C��2(�?E            �X@������������������������       �                     $@+       :                   �_@ą%�E�??            @V@,       -                    �?�IєX�?4             Q@������������������������       �        
             .@.       3                    \@�NW���?*            �J@/       2                    �L@�z�G��?             $@0       1                    @J@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @4       5                   `_@ qP��B�?"            �E@������������������������       �                     C@6       9                   �^@z�G�z�?             @7       8                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @;       @                   pb@���N8�?             5@<       ?                    �?�t����?	             1@=       >                    `@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     $@A       B                    �?      �?             @������������������������       �                     �?������������������������       �                     @D       O                    @Q@�t����?             1@E       H       
             �?z�G�z�?             .@F       G                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?I       J                    �?�8��8��?	             (@������������������������       �                      @K       L                   0r@ףp=
�?             $@������������������������       �                      @M       N                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @Q       R                   �X@��i#[�?             E@������������������������       �                      @S       Z                    �?��Q���?             D@T       Y                     P@�eP*L��?             &@U       X                    o@      �?              @V       W                   `_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @[       b                    �P@д>��C�?             =@\       ]       	          433�?HP�s��?             9@������������������������       �                     5@^       a                    �?      �?             @_       `                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?c       d                    �?      �?             @������������������������       �                     @������������������������       �                     �?f       �                    �?�=���?           �z@g       �                    �?:��0��?�            Pt@h       �       	          ���@����[��?2            �S@i       r       
             �?~X�<��?-             R@j       q                    �K@�q�q�?             (@k       p                    �E@      �?              @l       m                    \@      �?             @������������������������       �                      @n       o       	          @33�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @s       �       	             �?z�G�z�?"             N@t       }                   `\@V�a�� �?              M@u       z                   �c@      �?              @v       w                    �?z�G�z�?             @������������������������       �                     @x       y                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?{       |                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?~       �                   e@�:pΈ��?             I@       �                   �c@�X�<ݺ?             B@�       �                    �?��?^�k�?            �A@�       �                   0n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @@������������������������       �                     �?�       �                    �?X�Cc�?             ,@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                   �b@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �Q@���ʂ��?�            �n@�       �                   pf@�q�q�?             @�       �                    @G@�q�q�?             @������������������������       �                     �?�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	             @P�_��I�?�             n@�       �                    @L@�q3�M��?�             m@�       �       
             �?H��2�?s            @g@�       �       	          ����?     ��?             @@�       �                     F@      �?              @�       �                    `@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       
             �?      �?             8@�       �                   `]@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    @I@�}�+r��?             3@������������������������       �        	             (@�       �       	          033�?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    �J@�䞠�l�?]            @c@������������������������       �        H            �]@�       �                    �?��?^�k�?            �A@������������������������       �                     .@�       �                    @K@P���Q�?             4@�       �                   Hp@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     "@�       �       
             �?8����?             G@�       �                    @N@�q�q�?	             (@�       �       	          833�?�����H�?             "@������������������������       �                     @�       �                   `b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �^@@�0�!��?             A@������������������������       �                     "@�       �                    �?�+e�X�?             9@������������������������       �                     "@�       �                   `c@      �?
             0@�       �                     @"pc�
�?             &@�       �       	          @33�?z�G�z�?             $@������������������������       �                     @�       �                   p`@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    b@z�G�z�?             @������������������������       �                     @�       �                    e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �p@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                   �b@:ɨ��?<            �X@�       �                   �Z@b�h�d.�?)            �Q@������������������������       �                     @�       �                    f@�[|x��?&            �O@�       �                    �?P���Q�?$             N@�       �                   m@؇���X�?	             ,@������������������������       �                      @������������������������       �                     (@�       �       
             �?��<b�ƥ?             G@������������������������       �                     B@�       �       	             @ףp=
�?             $@�       �                   a@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �g@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    `@����"�?             =@�       �       	             �?      �?              @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @b@����X�?             5@�       �                   �q@     ��?	             0@�       �       
             �?�r����?             .@������������������������       �                     @�       �                    �?z�G�z�?             $@�       �                    a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �O@���Q��?             @������������������������       �                     @������������������������       �                      @�                          �^@� ��1�?}            �i@�       �                   @e@�U�:��?$            �M@�       �                    �? 7���B�?!             K@������������������������       �                    �F@�       �                    Z@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�       �       	          ����?���Q��?             @������������������������       �                      @�       �                    �H@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         �?f�Sa6T�?Y            @b@            
             �?���M�?8            @V@                        Pz@ ��PUp�?/            �Q@������������������������       �        .            �Q@������������������������       �                     �?                         �K@�E��ӭ�?	             2@                          F@X�<ݚ�?             "@������������������������       �                     @	      
                  @[@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@                        �o@6C�z��?!            �L@                        �`@p�ݯ��?             C@������������������������       �                     &@                        �O@�����H�?             ;@            	             �?      �?             @������������������������       �                      @������������������������       �                      @            	          ����?�nkK�?             7@                        ``@r�q��?             @������������������������       �                     @            
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     1@                        Pc@�d�����?             3@������������������������       �                     &@            	          033�?      �?              @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�B�       pz@     �~@     �w@     �t@     @U@     �i@      .@     �T@      *@      &@      @              @      &@      @      &@              $@      @      �?       @              �?      �?              �?      �?              @               @     �Q@      �?              �?     �Q@             �J@      �?      2@      �?      @              @      �?                      .@     �Q@     �^@      ;@      @      5@       @      4@              �?       @      �?                       @      @      @              @      @      �?       @      �?              �?       @              @             �E@     �\@      ,@     �Y@      "@     �V@              $@      "@      T@      @      P@              .@      @     �H@      @      @      @       @               @      @                      @      �?      E@              C@      �?      @      �?       @               @      �?                       @      @      0@       @      .@       @      @       @                      @              $@      @      �?              �?      @              @      (@      @      (@       @      �?       @                      �?      �?      &@               @      �?      "@               @      �?      �?      �?                      �?       @              =@      *@               @      =@      &@      @      @       @      @       @      �?       @                      �?              @      @              8@      @      7@       @      5@               @       @      �?       @               @      �?              �?              �?      @              @      �?             �r@     �_@     �p@     �L@     �J@      9@     �J@      3@      @      @      �?      @      �?      @               @      �?      �?              �?      �?                      @      @              H@      (@      G@      (@      @      @      �?      @              @      �?      �?              �?      �?               @      �?       @                      �?     �E@      @      A@       @      A@      �?       @      �?       @                      �?      @@                      �?      "@      @       @       @               @       @              @      @      @                      @       @                      @     �j@      @@       @      @       @      �?      �?              �?      �?              �?      �?                      @     �j@      <@     @j@      6@     @f@       @      9@      @      @      @      �?      @              @      �?              @              5@      @      @       @               @      @              2@      �?      (@              @      �?      @                      �?      c@      �?     �]@              A@      �?      .@              3@      �?      $@      �?      $@                      �?      "@              @@      ,@      @       @      �?       @              @      �?       @      �?                       @      @              <@      @      "@              3@      @      "@              $@      @      "@       @       @       @      @              @       @               @      @              �?              �?      @              @      �?      �?              �?      �?              @      @              @      @              >@     @Q@      (@      M@      @              @      M@      @     �L@       @      (@       @                      (@      �?     �F@              B@      �?      "@      �?      @      �?                      @              @       @      �?       @                      �?      2@      &@      @      @      �?      @              @      �?               @      �?              �?       @              .@      @      *@      @      *@       @      @               @       @       @       @       @                       @      @                      �?       @      @              @       @              D@     �d@      @      K@       @      J@             �F@       @      @       @                      @      @       @       @              �?       @      �?                       @     �A@     �[@      @     �T@      �?     �Q@             �Q@      �?              @      *@      @      @              @      @      �?              �?      @                      "@      =@      <@      8@      ,@              &@      8@      @       @       @               @       @              6@      �?      @      �?      @              �?      �?              �?      �?              1@              @      ,@              &@      @      @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ!�oZhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKۅ�h~�B�/         �       
             �?\r��ۖ�?K           ��@                          0b@\|/��j�?O           ��@       
                    �J@�z�N��?Q            ``@                          �a@`Ӹ����?            �F@������������������������       �                    �D@       	                    �?      �?             @                          �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?              	          033�?��f�{��?4            �U@������������������������       �        $             N@                           �? ��WV�?             :@������������������������       �        	             2@                          �]@      �?              @������������������������       �                     @              	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @       I                    �?Pw^�$C�?�            �x@       B                    �?Ȱi�o��?�            Pp@       )                    �?\-��p�?�            `i@              	          ����?�p ��?            �D@                           �?�θ�?             *@������������������������       �                      @              	            �?���Q��?             @������������������������       �                     @������������������������       �                      @       "                    �?X�Cc�?             <@       !                    �?���Q��?             $@                           �t@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @#       (                   �a@�<ݚ�?             2@$       '                    �J@      �?              @%       &                    �G@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     $@*       -                   �Z@H�!b	�?l            @d@+       ,                   �o@      �?             @������������������������       �                      @������������������������       �                      @.       /                    @J@(�5�f��?j            �c@������������������������       �        *            @P@0       ?                   �b@`Jj��?@            @W@1       6       	          ����?X;��?=            @V@2       3       	             �?8�Z$���?	             *@������������������������       �                     $@4       5                    j@�q�q�?             @������������������������       �                     �?������������������������       �                      @7       >                   `\@�"w����?4             S@8       9                   �[@���7�?             6@������������������������       �                     0@:       ;                    �?r�q��?             @������������������������       �                     @<       =                     M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        "             K@@       A                   �d@      �?             @������������������������       �                     @������������������������       �                     �?C       F                    �R@�8���?'             M@D       E                   �S@h�����?%             L@������������������������       �                      @������������������������       �        $             K@G       H                   p@      �?              @������������������������       �                     �?������������������������       �                     �?J       W                   a@�l�]�N�?T             a@K       R                    �?��2(&�?             F@L       M       	             �?      �?              @������������������������       �                     �?N       O                   �n@����X�?             @������������������������       �                     @P       Q                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?S       V                   �`@������?             B@T       U                   Pj@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     ;@X       q                   �`@\X��t�?7             W@Y       ^                    �?�-���?             I@Z       ]                   `c@�X�<ݺ?	             2@[       \                   @q@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@_       n       	          ���@      �?             @@`       k                    �?l��
I��?             ;@a       h       	             �?��<b���?             7@b       c                   �_@�t����?             1@������������������������       �                     *@d       g                    �?      �?             @e       f       	          833�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?i       j                    @      �?             @������������������������       �                     @������������������������       �                     @l       m       	            �?      �?             @������������������������       �                     @������������������������       �                     �?o       p       	             
@z�G�z�?             @������������������������       �                     @������������������������       �                     �?r       s       
             �?X�Cc�?             E@������������������������       �                     @t       �                   �d@      �?             B@u       |                    �?     ��?             @@v       w                   a@      �?              @������������������������       �                     @x       y                    �?z�G�z�?             @������������������������       �                     @z       {                    �?      �?              @������������������������       �                     �?������������������������       �                     �?}       ~                    �I@�8��8��?             8@������������������������       �                     ,@       �                    r@z�G�z�?             $@�       �                    �?�����H�?             "@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �N@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?���B���?�            `x@�       �                    �?x>ԛ/��?Q            �^@�       �                    @N@�n_Y�K�?A            �V@�       �                   @E@����?8            @S@�       �                    �?�n_Y�K�?
             *@�       �                    �?�q�q�?             @������������������������       �                     @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �L@և���X�?             @�       �                     E@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �a@     ��?.             P@������������������������       �                     7@�       �                   �_@v�2t5�?            �D@�       �                    �?�	j*D�?
             *@�       �                    �?      �?	             (@������������������������       �                      @�       �                   �n@ףp=
�?             $@������������������������       �                     @�       �                   0q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   �b@����X�?             <@�       �                    �?z�G�z�?             9@������������������������       �                     @�       �       	          `ff�?���N8�?             5@�       �                   �d@      �?             0@�       �                    `@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �                   @b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	          ����?����X�?	             ,@������������������������       �                     @�       �                     P@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �p@r֛w���?             ?@�       �       	          ����?HP�s��?             9@�       �                   ``@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �        	             .@������������������������       �                     @�       �                   0h@��	��j�?�            �p@�       �       	             @���}��?�            �p@�       �                    c@�.^J��?�            Pp@�       �                    c@����?�            �m@�       �       	            �?�θ�?             *@������������������������       �                     $@������������������������       �                     @�       �                   �^@���͡?�            @l@������������������������       �        <            �U@�       �                    _@��?^�k�?R            �a@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �i@`��(�?P            �`@�       �                    �?`Jj��?             ?@�       �                    @�8��8��?             8@������������������������       �                     6@������������������������       �                      @������������������������       �                     @������������������������       �        =             Z@�       �                    �?"pc�
�?             6@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@������������������������       �                     @�       �                    d@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       py@     �@      W@     @{@      @      `@       @     �E@             �D@       @       @       @      �?       @                      �?              �?      �?     @U@              N@      �?      9@              2@      �?      @              @      �?       @      �?                       @     @V@     @s@      ?@     �l@      <@     �e@      4@      5@      $@      @       @               @      @              @       @              $@      2@      @      @       @      @              @       @              @              @      ,@      @      @      @      �?              �?      @                      @              $@       @     @c@       @       @       @                       @      @      c@             @P@      @     �U@      @     �U@       @      &@              $@       @      �?              �?       @              �?     �R@      �?      5@              0@      �?      @              @      �?       @      �?                       @              K@      @      �?      @                      �?      @     �K@       @      K@       @                      K@      �?      �?              �?      �?              M@     �S@      @      C@      @      @              �?      @       @      @              �?       @               @      �?              �?     �A@      �?       @      �?                       @              ;@      J@      D@     �B@      *@      1@      �?      @      �?      @                      �?      $@              4@      (@      3@       @      2@      @      .@       @      *@               @       @       @      �?       @                      �?              �?      @      @              @      @              �?      @              @      �?              �?      @              @      �?              .@      ;@      @              "@      ;@      @      :@      @      @              @      @      �?      @              �?      �?      �?                      �?       @      6@              ,@       @       @      �?       @              @      �?       @              �?      �?      �?      �?                      �?      �?              @      �?              �?      @             �s@     �R@      P@      M@      L@     �A@      J@      9@      @       @       @      @              @       @      �?              �?       @              @      @      �?      @      �?                      @       @             �G@      1@      7@              8@      1@      @      "@      @      "@       @              �?      "@              @      �?       @      �?                       @      �?              4@       @      4@      @      @              0@      @      .@      �?      @      �?              �?      @              "@              �?      @              @      �?                      @      @      $@              @      @      @              @      @               @      7@       @      7@       @       @               @       @                      .@      @             `o@      1@     @o@      0@     @o@      &@      m@      @      $@      @      $@                      @     �k@      @     �U@              a@      @      @       @               @      @             �`@       @      =@       @      6@       @      6@                       @      @              Z@              2@      @      �?      @      �?                      @      1@                      @      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ[>tfhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK煔h~�B�2         �                    �?�6𿸴�?A           ��@       =                    �?@%�PWK�?a           ��@              
             �?��[�'�?�             i@                          �Q@P>�7���?G            @]@������������������������       �                      @                          `]@�LQ�1	�?F            �\@������������������������       �                    �C@                          (s@�=A�F�?.             S@	                          Pr@�jTM��?(            �N@
              	            �?F�t�K��?&            �L@������������������������       �                     9@                           �?     ��?             @@                          �^@r�q��?             8@������������������������       �                     @              	          ����?�����?             3@������������������������       �                     @              	          ����?�r����?             .@                          pm@�q�q�?             @                           �I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                      @������������������������       �                     @������������������������       �                     .@       $                   @E@�P�����?9             U@       #       	             �?؇���X�?             ,@       "                    �?      �?              @                          �X@      �?             @������������������������       �                     �?        !                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @%       <       	          ����?z��R[�?.            �Q@&       /                    �?��f/w�?(            �N@'       .                   Xv@�q�q�?	             (@(       -       	          @33�?z�G�z�?             $@)       ,                   �q@      �?              @*       +                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                      @0       1                   �k@ i���t�?            �H@������������������������       �                     8@2       ;                   �m@z�G�z�?             9@3       4                    �?�n_Y�K�?             *@������������������������       �                      @5       6                   �b@�eP*L��?             &@������������������������       �                     @7       :                   �l@r�q��?             @8       9                    �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                     "@>       M                   �O@�)l�o��?�            �v@?       L                    �?���@M^�?             ?@@       C                    �?�eP*L��?             6@A       B       	          ����?؇���X�?             @������������������������       �                     �?������������������������       �                     @D       K                    @���Q��?             .@E       F       	          �������
ц��?             *@������������������������       �                     @G       H                     P@�z�G��?             $@������������������������       �                     @I       J                   `]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@N       {       
             �?4�{Y���?�            �t@O       Z                    �?�W*��?7            @X@P       Q                   `Z@R���Q�?             4@������������������������       �                     �?R       S                   Pc@�KM�]�?             3@������������������������       �                     ,@T       U                   �`@���Q��?             @������������������������       �                      @V       Y                    �?�q�q�?             @W       X       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?[       `                   �k@*-ڋ�p�?)            @S@\       ]                   `g@r�q��?
             8@������������������������       �                      @^       _                    @�C��2(�?             6@������������������������       �                     4@������������������������       �                      @a       r                   �o@�F�j��?            �J@b       i       	            �?�+e�X�?             9@c       d       
             �?���Q��?             @������������������������       �                     �?e       f                    �O@      �?             @������������������������       �                      @g       h                   pm@      �?              @������������������������       �                     �?������������������������       �                     �?j       m                   �b@R���Q�?
             4@k       l                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?n       q                    �?�����H�?             2@o       p       
             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     *@s       z                   f@      �?             <@t       u                    �?�J�4�?             9@������������������������       �                     @v       w                    �J@���y4F�?             3@������������������������       �                     @x       y       
             �?�	j*D�?             *@������������������������       �                     @������������������������       �                     "@������������������������       �                     @|       �                    �?p�y�&z�?�            `m@}       �                   @c@������?            �B@~                          �`@      �?
             (@������������������������       �                     @�       �                    �?���Q��?             @�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       	          @33�?`2U0*��?             9@�       �                    �?�IєX�?             1@�       �                   �g@      �?              @������������������������       �                     @�       �                   pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                      @�       �                   @[@`�LVXz�?{            �h@�       �                    �?�<ݚ�?             "@������������������������       �                     @�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        u            �g@�       �       	          ����?p/3�d��?�             v@�       �                   �Y@�{ /h��?2            �S@�       �                    �?�}�+r��?             3@������������������������       �        	             *@�       �                    ^@r�q��?             @������������������������       �                     @�       �                    �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   Pd@�ݜ����?&            �M@�       �                    �?���3L�?#             K@�       �                   pb@�q�q�?             (@�       �                     N@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	          833�?X�Cc�?             E@�       �                   pq@�������?             A@�       �       
             �?8^s]e�?             =@������������������������       �                     1@�       �                    �?      �?             (@�       �                   �o@      �?              @������������������������       �                     @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     P@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   `^@      �?              @������������������������       �                     �?�       �                   �^@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?<���|��?�            @q@�       �                    �?      �?             <@�       �                   h@�q�q�?             5@�       �                    V@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                    �?      �?             0@�       �                    @I@ףp=
�?	             $@�       �                    �H@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	             �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    @G@��b�=�?�             o@�       �                    �C@"pc�
�?             6@������������������������       �                     @�       �                   �d@      �?             0@�       �                    \@؇���X�?
             ,@������������������������       �                      @������������������������       �        	             (@������������������������       �                      @�       �                    �?���=��?�            @l@�       �                    V@�X-:oȤ?v             h@������������������������       �                     @�       �       
             �?@_�M�q�?u            �g@�       �       	          033�?@�����?h             e@������������������������       �        /             S@�       �                   �b@�L��ȕ?9            @W@������������������������       �        4            �T@�       �                   �a@ףp=
�?             $@�       �       
             �?z�G�z�?             @������������������������       �                     �?�       �                     P@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     5@�       �                   �`@�'�`d�?            �@@�       �       
             �? �q�q�?             8@������������������������       �                     7@������������������������       �                     �?�       �                   `b@�q�q�?             "@������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp       �y@     p@     �v@      i@      S@     @_@      1@      Y@       @              .@      Y@             �C@      .@     �N@      .@      G@      &@      G@              9@      &@      5@      &@      *@      @              @      *@      @               @      *@       @      @       @      �?              �?       @                      @              "@               @      @                      .@     �M@      9@       @      (@       @      @       @       @              �?       @      �?              �?       @                      @              @     �L@      *@      H@      *@      @       @       @       @       @      @       @      �?              �?       @                      @               @       @              F@      @      8@              4@      @       @      @       @              @      @      @              �?      @      �?      �?              �?      �?                      @      (@              "@              r@     �R@      (@      3@      (@      $@      @      �?              �?      @              @      "@      @      @      @              @      @              @      @      �?      @                      �?               @              "@     @q@      L@     �G@      I@      1@      @              �?      1@       @      ,@              @       @       @              �?       @      �?      �?      �?                      �?              �?      >@     �G@      @      4@       @               @      4@              4@       @              :@      ;@      3@      @       @      @      �?              �?      @               @      �?      �?      �?                      �?      1@      @      �?      �?      �?                      �?      0@       @      @       @               @      @              *@              @      5@      @      5@              @      @      .@              @      @      "@      @                      "@      @             �l@      @     �@@      @      "@      @      @               @      @       @      �?              �?       @                       @      8@      �?      0@      �?      @      �?      @              �?      �?      �?                      �?      "@               @             �h@       @      @       @      @              �?       @               @      �?             �g@             �I@     �r@      =@     �H@      �?      2@              *@      �?      @              @      �?       @      �?                       @      <@      ?@      7@      ?@       @      @       @      @              @       @              @              .@      ;@      "@      9@      "@      4@              1@      "@      @      @      �?      @              �?      �?              �?      �?               @       @       @                       @              @      @       @              �?      @      �?      @                      �?      @              6@     �o@      @      5@      @      ,@      @       @               @      @              @      (@      �?      "@      �?      @              @      �?                      @      @      @      @                      @              @      .@      m@      @      2@              @      @      (@       @      (@       @                      (@       @              &@     �j@      @     �g@      @              �?     �g@      �?      e@              S@      �?      W@             �T@      �?      "@      �?      @              �?      �?      @      �?                      @              @              5@      @      :@      �?      7@              7@      �?              @      @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�BX7         V                   a@������?R           ��@              	             �?��b��a�?           �z@                           �?�G�z��?g             d@       	                   �h@     ��?             @@              	          @33�?      �?             $@                           �K@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @
                           �K@���7�?             6@������������������������       �                     .@              
             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @              
             �?     x�?S             `@              	          ����?�}#���?6            �T@                           �D@ ��PUp�?.            �Q@������������������������       �                     �?������������������������       �        -            �Q@                          �[@      �?             (@              
             �?�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @                           �M@�r����?            �F@              	             �?��?^�k�?            �A@������������������������       �                     A@������������������������       �                     �?                           �?      �?             $@������������������������       �                     @������������������������       �                     @        1                    �?�����?�            �p@!       *                    �?�LQ�1	�?             7@"       %                   0l@�q�q�?             "@#       $                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?&       )                   �r@r�q��?             @'       (                   @q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @+       0                    �?؇���X�?	             ,@,       -                    k@�q�q�?             @������������������������       �                      @.       /                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @2       S                    @0 �����?�            @n@3       P                    �R@@Ix�<��?�            �m@4       K       
             �?xsG��?�             m@5       @                   `_@p� V�?�            �i@6       7                    �?�"w����?e             c@������������������������       �        G            �Z@8       ?                   �`@`Ӹ����?            �F@9       :                   �X@z�G�z�?             $@������������������������       �                     �?;       >       
             �?�����H�?             "@<       =                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                    �A@A       F                     E@ 7���B�?"             K@B       C                    b@؇���X�?             @������������������������       �                     @D       E                    �C@�q�q�?             @������������������������       �                      @������������������������       �                     �?G       J                    \@`Ql�R�?            �G@H       I       	          033@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     F@L       M                   �_@������?             ;@������������������������       �                     3@N       O                     P@      �?              @������������������������       �                     @������������������������       �                     �?Q       R       	             @      �?             @������������������������       �                      @������������������������       �                      @T       U                    �?���Q��?             @������������������������       �                     @������������������������       �                      @W       �                    �?p�NO���??           �~@X       �       
             �?nj���X�?�             x@Y       r                    @L@�p�o�?�?L            �[@Z       a                    �?�)�8��?0             Q@[       `                    �H@�IєX�?             1@\       _                   �_@z�G�z�?             @]       ^                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@b       q                   �f@j���� �?$            �I@c       d                    �?�LQ�1	�?!             G@������������������������       �                     *@e       j                    �?�'�=z��?            �@@f       g                     H@     ��?	             0@������������������������       �                     &@h       i       	          ����?���Q��?             @������������������������       �                     @������������������������       �                      @k       p                    �K@@�0�!��?             1@l       o                   �a@      �?             0@m       n                   @g@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             &@������������������������       �                     �?������������������������       �                     @s       �                   �e@>��C��?            �E@t       u       
             �?d}h���?             E@������������������������       �                     $@v       �                   �b@     ��?             @@w       �                    b@��H�}�?             9@x       y                   b@8����?             7@������������������������       �                     @z       �                    �N@j���� �?             1@{       �                    �?"pc�
�?             &@|       }                   �b@�<ݚ�?             "@������������������������       �                     �?~                           �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?r�q��?             @������������������������       �                     @�       �                   Pn@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �       	          `ff @�;�a
=�?�            0q@�       �                    �? �N����?�            �p@�       �                    �?� ���?(            @P@�       �                    b@θ	j*�?"             J@�       �                   �a@��Sݭg�?            �C@������������������������       �        	             &@�       �                   �c@X�Cc�?             <@�       �       	          @33�?�eP*L��?             &@�       �                    �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �s@������?             1@�       �                    �?$�q-�?
             *@������������������������       �                     "@�       �                   d@      �?             @�       �                   Pm@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �L@��
ц��?             *@�       �                     E@����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     �?�       �                   `Y@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �a@$�q-�?             *@�       �       	          hff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�       �                   �t@г�wY;�?            �i@�       �                   `i@@�E�x�?y            �h@������������������������       �        #            �N@�       �       	          ����?@A��q�?V            �`@�       �                   @[@P�c0"�?F            @Z@�       �                     H@r�q��?             @�       �                    @D@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?`�LVXz�?@            �X@�       �                   `b@�X�<ݺ?
             2@������������������������       �                     0@�       �                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        6            @T@�       �                   �a@��S�ۿ?             >@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    j@h�����?             <@�       �                     I@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     8@�       �                    �?      �?              @�       �                   u@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?"�a�5M�?H            �Z@�       �                   pl@�{ /h��?7            �S@�       �                    �?�c�Α�?             =@�       �                   `e@r�q��?             8@�       �                    c@�LQ�1	�?             7@�       �       
             �?�θ�?
             *@�       �                    �?"pc�
�?             &@������������������������       �                     @�       �                    �H@      �?              @������������������������       �                      @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     �?�       �                    e@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	            �?ZՏ�m|�?"            �H@�       �                   pb@��
ц��?             *@������������������������       �                     @�       �                   `c@���Q��?             $@������������������������       �                     @�       �                   `d@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                   �[@�X�<ݺ?             B@�       �                    �?؇���X�?             @������������������������       �                     @�       �                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    q@XB���?             =@������������������������       �                     .@�       �       	          ����?@4և���?             ,@������������������������       �                     "@�       �                    c@z�G�z�?             @������������������������       �                     @�       �                    �J@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	             �?\-��p�?             =@�       �                    �I@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     6@�t�b��     h�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@      X@     �t@      R@      V@      :@      @      @      @       @      @       @                      @      @              5@      �?      .@              @      �?              �?      @              G@     �T@      @      S@      �?     �Q@      �?                     �Q@      @      @      @      @      @                      @      @             �C@      @      A@      �?      A@                      �?      @      @              @      @              8@      n@       @      .@      @      @      �?       @               @      �?              @      �?       @      �?       @                      �?      @               @      (@       @      @               @       @       @       @                       @               @      0@     @l@      *@      l@      &@     �k@      @     @i@       @     �b@             �Z@       @     �E@       @       @      �?              �?       @      �?       @               @      �?                      @             �A@       @      J@      �?      @              @      �?       @               @      �?              �?      G@      �?       @      �?                       @              F@      @      4@              3@      @      �?      @                      �?       @       @       @                       @      @       @      @                       @     �s@     `f@     �q@     @Z@     �G@      P@     �B@      ?@      0@      �?      @      �?      �?      �?      �?                      �?      @              (@              5@      >@      0@      >@              *@      0@      1@      *@      @      &@               @      @              @       @              @      ,@       @      ,@       @      @       @                      @              &@      �?              @              $@     �@@      "@     �@@              $@      "@      7@      "@      0@      @      0@              @      @      $@       @      "@       @      @      �?              �?      @              @      �?                       @      @      �?      @               @      �?       @                      �?       @                      @      �?             @m@     �D@     @m@     �A@      B@      =@     �A@      1@      =@      $@      &@              2@      $@      @      @      @       @               @      @                      @      *@      @      (@      �?      "@              @      �?      �?      �?              �?      �?               @              �?      @              @      �?              @      @      @       @               @      @              �?      @              �?      �?      @      �?                      @      �?      (@      �?      �?      �?                      �?              &@     �h@      @      h@      @     �N@             ``@      @     �Y@       @      @      �?       @      �?       @                      �?      @             �X@      �?      1@      �?      0@              �?      �?              �?      �?             @T@              <@       @      �?      �?              �?      �?              ;@      �?      @      �?      @                      �?      8@              @       @      @       @               @      @               @                      @     �@@     �R@      =@     �H@      5@       @      4@      @      4@      @      $@      @      "@       @      @              @       @               @      @              �?      �?              �?      �?              $@                      �?      �?      @              @      �?               @     �D@      @      @              @      @      @      @               @      @              @       @               @      A@      �?      @              @      �?      �?      �?                      �?      �?      <@              .@      �?      *@              "@      �?      @              @      �?      �?              �?      �?              @      9@      @      @              @      @                      6@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJy-ahG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKׅ�h~�B/         ~       
             �?��t�?J           ��@       K                    �?fP*L��?U           ��@                           �F@,˫�5�?�            �h@                           �?D^��#��?            �D@       
                    ]@�<ݚ�?
             2@                          �Z@z�G�z�?             @������������������������       �                      @       	                    �D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@                          �[@��<b���?             7@������������������������       �                     @                           @ףp=
�?             4@                          @^@�}�+r��?             3@                          �o@      �?              @������������������������       �                     @                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@������������������������       �                     �?       *                    �?������?o            �c@                            L@��S���?            �F@              	          ����?$�q-�?             *@������������������������       �                     (@������������������������       �                     �?       '                    @     ��?             @@                            @P@d}h���?             <@                          �Z@�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@!       &                   �b@      �?             $@"       #                    �?����X�?             @������������������������       �                      @$       %                   @L@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @(       )                   `\@      �?             @������������������������       �                     �?������������������������       �                     @+       .       	          833�?�SM:$�?P            @\@,       -       
             �?@��8��?!             H@������������������������       �                     �?������������������������       �                     �G@/       B                   �`@��&����?/            @P@0       1       	             �?`՟�G��?             ?@������������������������       �                     @2       5                    �?��>4և�?             <@3       4                   `_@؇���X�?
             ,@������������������������       �                     (@������������������������       �                      @6       7       
             �?X�Cc�?             ,@������������������������       �                     �?8       ?                   �n@�	j*D�?
             *@9       >                    e@z�G�z�?             $@:       =                   �W@�����H�?             "@;       <                    �M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?@       A                   Xr@�q�q�?             @������������������������       �                      @������������������������       �                     �?C       J                    �?l��\��?             A@D       E                    �I@�LQ�1	�?             7@������������������������       �                      @F       I       	          ����?z�G�z�?
             .@G       H                    X@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                     &@L       }       	          `ff @H�E�@��?�            �t@M       Z                   �[@�C��2(�?�            �o@N       S                   `_@�q�q�?             8@O       P                    �?ףp=
�?             $@������������������������       �                     @Q       R       	          `ff�?      �?             @������������������������       �                     @������������������������       �                     �?T       U                    �?X�Cc�?	             ,@������������������������       �                     @V       Y                    �?"pc�
�?             &@W       X                   �n@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @[       d                    �?����]j�?�            �l@\       a                    �?r�q��?             8@]       `       	          ����?ףp=
�?             4@^       _                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        
             ,@b       c                   �o@      �?             @������������������������       �                      @������������������������       �                      @e       z                   `f@��?ȿ}�?�            �i@f       w                    c@��*Td`�?            �h@g       v                    �R@@�.L3خ?{             h@h       u       	          ����?�X�T���?z            �g@i       j                    @L@�kb97�?4            @S@������������������������       �                     @@k       r                    �?�:�^���?            �F@l       q                   �X@�X�<ݺ?             B@m       n                    �?r�q��?             (@������������������������       �                      @o       p                   �W@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     8@s       t                    �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �        F            �\@������������������������       �                      @x       y                   `c@r�q��?             @������������������������       �                     �?������������������������       �                     @{       |                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        +             S@       �                    I@���B���?�            `x@�       �                    �?����X�?             E@�       �                    �?
;&����?             7@�       �                     E@     ��?	             0@������������������������       �                      @�       �                   @_@d}h���?             ,@������������������������       �                     @�       �                   �Y@      �?              @������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@�       �                    �L@X�
����?�            �u@�       �                    �?��S�ۿ?�            �p@�       �                   �a@��6}��?'            �N@�       �                    �?h�����?             <@�       �                    �I@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     3@�       �                    �?�eP*L��?            �@@�       �                   �_@`�Q��?             9@�       �                    �?���Q��?             $@������������������������       �                     @�       �                    �?؇���X�?             @�       �                   @^@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �b@�r����?	             .@������������������������       �                     *@������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                   @[@ �si�?�             j@�       �                   �l@��S�ۿ?             .@������������������������       �                     &@�       �                   @c@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �? �m�+�?y            @h@������������������������       �        (             P@�       �                    @L@��G^�C�?Q            @`@������������������������       �        O             `@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?$��m��?2            �S@�       �       	             �?��6}��?%            �N@�       �                    �N@D>�Q�?!             J@�       �                   pd@����X�?             <@�       �                   d@�ՙ/�?             5@�       �                    �?z�G�z�?             .@�       �                    _@      �?             @������������������������       �                     �?�       �                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�C��2(�?             &@�       �                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   0d@r�q��?             @������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     P@ �q�q�?             8@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                    �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@�       �                     Q@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    �?ҳ�wY;�?             1@�       �                   �q@�8��8��?	             (@������������������������       �                     $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp       �x@     8�@      U@     �{@     �N@     @a@      6@      3@      @      ,@      @      �?       @               @      �?              �?       @                      *@      2@      @              @      2@       @      2@      �?      @      �?      @               @      �?              �?       @              &@                      �?     �C@     �]@      5@      8@      (@      �?      (@                      �?      "@      7@      @      6@      �?      1@      �?                      1@      @      @       @      @               @       @      @       @                      @      @              @      �?              �?      @              2@     �W@      �?     �G@      �?                     �G@      1@      H@      ,@      1@      @              &@      1@       @      (@              (@       @              "@      @              �?      "@      @       @       @       @      �?       @      �?              �?       @              @                      �?      �?       @               @      �?              @      ?@      @      4@               @      @      (@      @      �?              �?      @                      &@              &@      7@      s@      7@     �l@      $@      ,@      �?      "@              @      �?      @              @      �?              "@      @              @      "@       @      @       @      @                       @      @              *@      k@      @      4@       @      2@       @      @              @       @                      ,@       @       @       @                       @      "@     �h@      @      h@      @     `g@      @     `g@      @     @R@              @@      @     �D@       @      A@       @      $@               @       @       @               @       @                      8@       @      @              @       @                     �\@       @              �?      @      �?                      @       @      @              @       @                      S@     �s@     �R@      (@      >@      (@      &@      @      &@       @              @      &@              @      @      @              @      @      �?      @                      �?      @                      3@     �r@     �F@     �o@      2@     �F@      0@      ;@      �?       @      �?              �?       @              3@              2@      .@      1@       @      @      @      @              �?      @      �?      @              @      �?                      �?      *@       @      *@                       @      �?      @      �?                      @     �i@       @      ,@      �?      &@              @      �?              �?      @              h@      �?      P@              `@      �?      `@              �?      �?              �?      �?             �I@      ;@     �F@      0@     �E@      "@      4@       @      *@       @      (@      @       @       @      �?              �?       @      �?                       @      $@      �?       @      �?              �?       @               @              �?      @              @      �?      �?              �?      �?              @              7@      �?      "@      �?      @               @      �?       @                      �?      ,@               @      @              @       @              @      &@      �?      &@              $@      �?      �?      �?                      �?      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJﴷ&hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�BX7         �       
             �?>���i��?^           ��@       %                    �?j��>��?Z           `�@                           �?��q7L��?;            �T@                          �V@ �o_��?$             I@������������������������       �                     @                          �p@�X����?              F@                           @M@� �	��?             9@       	                    �?ҳ�wY;�?             1@������������������������       �                     @
                           i@�eP*L��?             &@������������������������       �                     @              	             �?؇���X�?             @                          �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @                           �?�S����?             3@                          �x@��S�ۿ?             .@������������������������       �                     &@              	          ����?      �?             @������������������������       �                     �?������������������������       �                     @                           �?      �?             @������������������������       �                     �?              	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       $                    �?�'�`d�?            �@@       #                   `c@@4և���?             <@       "       	          ����? 7���B�?             ;@        !                   �e@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@������������������������       �                     �?������������������������       �                     @&       �       	          ���@`�C�h��?           �{@'       :                    e@4?,R��?�            �v@(       7                    �Q@�d���Ҹ?U             a@)       0       	          033�?5�wAd�?S            �`@*       +                    �?`�LVXz�?<            �X@������������������������       �        0             S@,       /                   `X@�nkK�?             7@-       .                    V@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             3@1       2                   �]@(N:!���?            �A@������������������������       �                     3@3       4                   �^@      �?
             0@������������������������       �                     "@5       6                    �?և���X�?             @������������������������       �                     @������������������������       �                     @8       9                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?;       F       
             �?h�!��?�            �k@<       A       	          ����?      �?             4@=       >                    d@      �?              @������������������������       �                     @?       @                   e@      �?              @������������������������       �                     �?������������������������       �                     �?B       C                    �?      �?	             (@������������������������       �                     @D       E                     O@���Q��?             @������������������������       �                      @������������������������       �                     @G       r                   pn@J'���l�?�            `i@H       S                   `_@�le����?G            �Z@I       L                   @\@���U�?$            �L@J       K                    �?      �?              @������������������������       �                     �?������������������������       �                     �?M       N                    �? �Jj�G�?"            �K@������������������������       �                    �C@O       R                    �?      �?             0@P       Q                   `Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@T       ]                   �]@�q�����?#             I@U       Z                   �m@8�Z$���?             *@V       Y                    �?�C��2(�?             &@W       X                    b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @[       \                    �?      �?              @������������������������       �                     �?������������������������       �                     �?^       q                    �?^H���+�?            �B@_       l                    �?П[;U��?             =@`       e                    �?b�2�tk�?             2@a       d                    �?���Q��?             @b       c                   0a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @f       k                    m@�n_Y�K�?             *@g       j       	          ����?z�G�z�?             $@h       i                   @`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @m       n                   Pf@"pc�
�?
             &@������������������������       �                     �?o       p                   `b@ףp=
�?	             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                      @s       �                   @^@�8��8N�?B             X@t       {                   �r@      �?             @@u       z                   0p@ ��WV�?             :@v       w                   �a@r�q��?             @������������������������       �                     @x       y                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@|       }                   `]@      �?             @������������������������       �                      @~                           �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   q@     �?+             P@������������������������       �                     9@�       �                   �e@$�q-�?            �C@�       �                    �?�?�|�?            �B@������������������������       �                     "@�       �                   �b@h�����?             <@������������������������       �                     ;@������������������������       �                     �?������������������������       �                      @�       �                   �i@F|/ߨ�?3            @T@������������������������       �                     B@�       �                    j@`Ӹ����?            �F@������������������������       �                     �?�       �                    �?`���i��?             F@������������������������       �                     B@�       �       
             �?      �?              @������������������������       �                      @�       �                   �`@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   @E@���5��?           �x@�       �                   P`@�q����?            �J@�       �                    �?�r����?             >@������������������������       �                     4@�       �                   pf@���Q��?             $@�       �       	          �ff�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �`@
;&����?             7@������������������������       �                     @�       �                   �a@b�2�tk�?	             2@�       �       	          ����?���!pc�?             &@�       �                    �?և���X�?             @�       �                    [@�q�q�?             @������������������������       �                      @�       �                   �]@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?և���X�?             @�       �       	          ���@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?�H�KY�?�            Pu@�       �       	          033@p���?�            �r@�       �                    �?˒�#�?�            �r@�       �                    q@8��8���?"             H@�       �                    �?�8��8��?             B@�       �                    �K@�S����?             3@�       �                   i@��S�ۿ?	             .@�       �                     B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@�       �                   �b@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     1@�       �                   �r@�q�q�?
             (@������������������������       �                     @�       �                    t@�����H�?             "@�       �                   �s@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?�a�n`�?�             o@������������������������       �        8            �W@�       �                   �_@���7�?k            @c@�       �                   �^@85�}C�?,            �N@�       �                    ]@ ��WV�?&             J@�       �                   c@ףp=
�?             4@�       �                   �[@z�G�z�?             $@�       �                    j@�����H�?             "@������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   �n@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     @@�       �                    �?�q�q�?             "@������������������������       �                     �?�       �                    _@      �?              @�       �                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �c@����D��??            @W@������������������������       �        (            �K@�       �                   xt@�}�+r��?             C@�       �                   Pd@��?^�k�?            �A@�       �                     L@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     9@�       �                   Xw@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �M@X��ʑ��?!            �E@�       �       	          033�?��}*_��?             ;@�       �                    �?��+7��?             7@�       �                   @d@��
ц��?	             *@�       �                    �?�q�q�?             "@�       �                    n@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   `a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �        
             $@������������������������       �                     @�       �                   Pp@      �?             0@������������������������       �                      @�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@      W@      {@      D@     �E@      ,@      B@              @      ,@      >@      &@      ,@      &@      @      @              @      @      @              �?      @      �?      �?      �?                      �?              @               @      @      0@      �?      ,@              &@      �?      @      �?                      @       @       @              �?       @      �?       @                      �?      :@      @      :@       @      :@      �?      @      �?      @                      �?      3@                      �?              @      J@     Px@      I@     `s@      @     @`@      @      `@      �?     �X@              S@      �?      6@      �?      @              @      �?                      3@      @      ?@              3@      @      (@              "@      @      @              @      @               @      �?       @                      �?     �E@     �f@      $@      $@      @      �?      @              �?      �?              �?      �?              @      "@              @      @       @               @      @             �@@     @e@      :@     @T@       @     �K@      �?      �?              �?      �?              �?      K@             �C@      �?      .@      �?      @      �?                      @              "@      8@      :@      &@       @      $@      �?      @      �?      @                      �?      @              �?      �?              �?      �?              *@      8@      *@      0@      &@      @      @       @      �?       @      �?                       @       @               @      @       @       @      �?       @               @      �?              @                      @       @      "@      �?              �?      "@              "@      �?                       @      @     @V@      @      <@      �?      9@      �?      @              @      �?      �?      �?                      �?              4@      @      @       @              �?      @      �?                      @      @     �N@              9@      @      B@      �?      B@              "@      �?      ;@              ;@      �?               @               @     �S@              B@       @     �E@      �?              �?     �E@              B@      �?      @               @      �?      @      �?                      @     �s@     �R@      0@     �B@      @      :@              4@      @      @      @      �?      @                      �?              @      (@      &@      @              @      &@      @       @      @      @       @      @               @       @       @       @                       @      �?                      @      @      @       @      @       @                      @       @             �r@      C@     �q@      0@     �q@      ,@     �D@      @     �@@      @      0@      @      ,@      �?      �?      �?      �?                      �?      *@               @       @      �?              �?       @      �?                       @      1@               @      @              @       @      �?      @      �?      @                      �?      @              n@      @     �W@             `b@      @      L@      @      I@       @      2@       @       @       @       @      �?      @              @      �?       @               @      �?              �?       @                      �?      $@              @@              @      @              �?      @       @      �?       @               @      �?              @             �V@       @     �K@              B@       @      A@      �?      "@      �?      "@                      �?      9@               @      �?              �?       @                       @      5@      6@      1@      $@      1@      @      @      @      @      @      �?      @      �?                      @       @       @               @       @              @              $@                      @      @      (@               @      @      @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�pD=hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�:         �                    �?\r��ۖ�?K           ��@       Y       
             �?*��r��?6           �~@       T                    �Q@��}�?�            �w@                           �?���UC5�?�            Pw@                           �J@^(��I�?#            �K@                           �D@�G�z��?             4@������������������������       �                     @       	                   �k@X�Cc�?
             ,@������������������������       �                     @
                           @I@"pc�
�?             &@������������������������       �                      @                            J@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?؇���X�?            �A@                           �?����X�?             ,@                           @O@      �?              @                           �N@�q�q�?             @������������������������       �                     �?                          �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @              	          033�?      �?             @������������������������       �                     @������������������������       �                     @                           �?���N8�?             5@������������������������       �                     0@              	          hff�?z�G�z�?             @������������������������       �                     �?������������������������       �                     @        -                    �?x��-�?�            �s@!       &                   pr@ܷ��?��?3            �U@"       #       	          833�?`<)�+�?,            @S@������������������������       �                     I@$       %       	          033�?�����H�?             ;@������������������������       �                     @������������������������       �                     8@'       *       
             �?���Q��?             $@(       )                    �?      �?             @������������������������       �                      @������������������������       �                      @+       ,                   @_@�q�q�?             @������������������������       �                     @������������������������       �                      @.       O                    c@���N8�?�            �l@/       6       	          ����?`2U0*��?�             l@0       1       	          833�?$G$n��?            �B@������������������������       �                     =@2       3                   �Y@      �?              @������������������������       �                      @4       5                   @_@r�q��?             @������������������������       �                     @������������������������       �                     �?7       F                   pa@`Ql�R�?y            �g@8       =       	          033@�e���@�?e            @c@9       <                   0i@ 
�V�?V            �`@:       ;                   h@ �.�?Ƞ?$             N@������������������������       �        #            �M@������������������������       �                     �?������������������������       �        2            �R@>       ?                    �?P���Q�?             4@������������������������       �        
             (@@       E       	             @      �?              @A       D                    ]@z�G�z�?             @B       C                     M@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @G       N                   �a@�IєX�?             A@H       I                    �?r�q��?             (@������������������������       �                     @J       K       
             �?      �?              @������������������������       �                      @L       M                    �H@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     6@P       Q                    q@�q�q�?             @������������������������       �                     @R       S                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?U       V                   `g@      �?             @������������������������       �                     �?W       X                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?Z       e                   �c@��"Ӗ��?H            @]@[       d                   �`@z�G�z�?            �A@\       c                   �_@p�ݯ��?             3@]       ^                   �_@z�G�z�?	             .@������������������������       �                      @_       b                    �N@և���X�?             @`       a       	             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        	             0@f       s                    �?��p �?4            �T@g       r                   �v@��}*_��?             ;@h       i                   �Y@�q�q�?             8@������������������������       �                     @j       k                     G@��s����?             5@������������������������       �                     @l       q       	          @33�?      �?             0@m       n                    `@      �?              @������������������������       �                      @o       p                   pe@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @t                           �?t�6Z���?$            �K@u       z                    @L@@4և���?             E@v       y                    �D@������?             B@w       x                    @C@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     =@{       ~                    �O@�q�q�?             @|       }                   @g@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   b@�n_Y�K�?	             *@�       �                   �[@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             @�       �                   pd@���Q��?             @�       �                   Hq@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �K@4S�t ��?           �z@�       �       
             �?8zw"׷�?�            @q@�       �                    @G@��.k���?*             Q@�       �                   �a@������?             >@�       �                   �[@����X�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   Pd@�LQ�1	�?             7@�       �                    �?�z�G��?             $@�       �                    c@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     *@�       �                    �?p�ݯ��?             C@�       �       	          ����?�q�q�?             (@������������������������       �                     @������������������������       �                      @�       �                    @J@�θ�?             :@�       �                   �m@���Q��?	             .@�       �       	             �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @�       �                   �`@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@�       �                    �?���%�?�             j@������������������������       �        -             Q@�       �       	             @h�����?W            �a@�       �                   c@��*����?V            `a@�       �                   @n@�>����?!             K@�       �       	          pff�?�(\����?             D@������������������������       �                    �B@�       �                    d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �n@d}h���?             ,@������������������������       �                     @������������������������       �                     &@������������������������       �        5            @U@������������������������       �                     �?�       �       
             �?��%��?g            �b@�       �                   �[@N�zv�?<             V@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @0,Tg��?9             U@�       �                   �b@@���?T�?-            �Q@�       �                   r@��mo*�?&            �M@�       �                   Pg@���y4F�?%            �L@�       �                    �?      �?
             0@�       �                    �L@؇���X�?             @�       �       	             �      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �                   @]@���� �?            �D@�       �                    �?      �?              @�       �                   �`@�q�q�?             @�       �       	          033�?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �       	          ����?�'�`d�?            �@@�       �       
             �?�����?             3@������������������������       �                     �?�       �       	          ����?�E��ӭ�?             2@�       �                   p@      �?              @������������������������       �                     @������������������������       �                     �?�       �                   �o@���Q��?             $@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �`@@4և���?	             ,@�       �                    @N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                      @�       �                   @]@�8��8��?             (@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                     M@��
ц��?             *@������������������������       �                      @�       �                    @O@�eP*L��?
             &@�       �       
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �k@�q�q�?             @������������������������       �                     �?�       �                     P@z�G�z�?             @������������������������       �                     @�       �                    p@      �?              @������������������������       �                     �?������������������������       �                     �?�             	          ����?��0u���?+             N@�       �       	          ����?�{��?��?(             K@�       �                    �?�c�Α�?             =@�       �                     R@`�Q��?             9@�       �                   �s@��+7��?             7@�       �                    c@R���Q�?             4@������������������������       �        
             .@�       �                    @N@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @                          �M@H%u��?             9@                        �p@�q�q�?             @                          M@�q�q�?             @                        �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        `Q@�}�+r��?             3@	      
      	          ����?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�B�       py@     �@      Y@     �x@      B@     Pu@      A@     0u@      ,@     �D@      "@      &@              @      "@      @              @      "@       @       @              �?       @               @      �?              @      >@      @      $@      �?      @      �?       @              �?      �?      �?      �?                      �?              @      @      @              @      @              �?      4@              0@      �?      @      �?                      @      4@     �r@      "@     �S@      @     �R@              I@      @      8@      @                      8@      @      @       @       @       @                       @      @       @      @                       @      &@     �k@      "@      k@      @      @@              =@      @      @               @      @      �?      @                      �?      @      g@       @      c@      �?     �`@      �?     �M@             �M@      �?                     �R@      �?      3@              (@      �?      @      �?      @      �?      @      �?                      @              �?              @       @      @@       @      $@              @       @      @               @       @      @       @                      @              6@       @      @              @       @      �?       @                      �?       @       @      �?              �?       @               @      �?              P@     �J@      @      <@      @      (@      @      (@               @      @      @      @      �?      @                      �?              @      @                      0@     �L@      9@      $@      1@      @      1@      @              @      1@              @      @      (@      @      @       @               @      @              @       @                       @      @             �G@       @     �C@      @     �A@      �?      @      �?      @                      �?      =@              @       @      �?       @      �?                       @      @               @      @      @      �?              �?      @               @      @       @      @      �?      @              @      �?              �?                      �?     0s@     @]@     �m@     �B@      B@      @@      6@       @       @      @              @       @      �?       @                      �?      4@      @      @      @       @      @       @                      @      @              *@              ,@      8@       @      @              @       @              @      4@      @      "@       @       @       @                       @      @      �?      @                      �?              &@     `i@      @      Q@             �`@      @     �`@      @      I@      @     �C@      �?     �B@               @      �?              �?       @              &@      @              @      &@             @U@                      �?      Q@      T@      9@     �O@      @      �?              �?      @              6@      O@      .@      L@      ,@     �F@      (@     �F@      �?      .@      �?      @      �?      �?              �?      �?                      @              "@      &@      >@      @      @      @       @       @       @               @       @               @                       @      @      :@      @      *@      �?              @      *@      �?      @              @      �?              @      @      @       @               @      @                      @      �?      *@      �?      @              @      �?                      "@       @              �?      &@      �?      @      �?                      @              @      @      @       @              @      @      �?      @      �?                      @      @       @              �?      @      �?      @              �?      �?      �?                      �?     �E@      1@     �E@      &@      5@       @      1@       @      1@      @      1@      @      .@               @      @              @       @                      @               @      @              6@      @      @       @      �?       @      �?      �?      �?                      �?              �?      @              2@      �?      @      �?      @                      �?      ,@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�XhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B(5         �                   �b@2���xA�?7           ��@       g       
             �?�E�p�?�           Ȅ@       `                    �Q@��p���?            }@                           �?Q9w2��?           `|@                          �`@��>4և�?!             L@       	       	          ����?`՟�G��?             ?@                           �N@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?
                           �O@������?             1@                           �J@؇���X�?             ,@                           �I@���Q��?             @                          �a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@                          `Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �I@z�G�z�?             9@              	             �?      �?              @������������������������       �                     @������������������������       �                     @                           `P@�IєX�?             1@������������������������       �        
             .@                          @\@      �?              @������������������������       �                     �?������������������������       �                     �?       S                    �?�h��$�?�            �x@       <                   `a@�1����?�            `p@        '       
             �?���a�\�?}            @i@!       &                   �U@r�q��?             8@"       %       	             �?�q�q�?             (@#       $                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     (@(       7       	          ���@ d���W�?p            @f@)       *                   �_@������?f            `d@������������������������       �        !            �J@+       6                   �p@h㱪��?E            �[@,       -                     E@ >�֕�?.            �Q@������������������������       �                      @.       5                   �[@г�wY;�?,             Q@/       4       	             �?�C��2(�?             6@0       3                    b@����X�?             @1       2                   �\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     .@������������������������       �                     G@������������������������       �                     D@8       9                    �?z�G�z�?
             .@������������������������       �                     $@:       ;                   p`@���Q��?             @������������������������       �                     @������������������������       �                      @=       R                   �b@���*�?$             N@>       G       	          ����?0,Tg��?             E@?       @                   �g@��
ц��?             *@������������������������       �                     @A       F                   �^@���Q��?             $@B       E                    �?z�G�z�?             @C       D                    @F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @H       M                    �?\-��p�?             =@I       L                   �j@���7�?             6@J       K                    b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             2@N       Q                    �N@և���X�?             @O       P       	          `ff @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �        
             2@T       ]                     Q@�����?K             a@U       Z                   Pz@@��A1ʞ?G            ``@V       W                    @�7�	|��?E             `@������������������������       �        B            @_@X       Y       	          `ff�?      �?             @������������������������       �                     @������������������������       �                     �?[       \                     L@      �?              @������������������������       �                     �?������������������������       �                     �?^       _       	          ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @a       b                    �?���Q��?             $@������������������������       �                     @c       d       	          033�?�q�q�?             @������������������������       �                      @e       f                    �?      �?             @������������������������       �                      @������������������������       �                      @h       �                    �?$@e����?�             i@i       �                   �_@6YE�t�?j            �d@j       w                   �e@     ��?$             P@k       l                    @H@��Q��?
             4@������������������������       �                      @m       v                    ^@�E��ӭ�?	             2@n       s                    �?      �?             $@o       r       	          ����?�q�q�?             @p       q                    �L@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @t       u                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @x                           @��2(&�?             F@y       z                    �?��(\���?             D@������������������������       �                     ?@{       ~                    �?�q�q�?             "@|       }                    o@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �K@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?(a��䛼?F            @Y@�       �       	          ����?"pc�
�?            �@@������������������������       �                     6@�       �                   �m@�eP*L��?             &@�       �                   �`@����X�?             @������������������������       �                     @�       �                   0k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �        .             Q@�       �                    �?b�2�tk�?             B@�       �                   @V@      �?              @������������������������       �                     �?������������������������       �                     @�       �                   �a@      �?             <@�       �       	          hff�?��Q��?             4@�       �                    �?���|���?             &@�       �                    �L@�<ݚ�?             "@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �                      @�       �                    @G@T<;="��?�            �o@�       �                   �[@8��8���?B             X@�       �                   @[@�eP*L��?
             &@�       �                    �?r�q��?             @������������������������       �                     @�       �                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     E@z�G�z�?             @������������������������       �                     @�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	             �?�̨�`<�?8            @U@�       �                   �c@�}�+r��?4             S@�       �                    �?�q�q�?             "@�       �       
             �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   q@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   hq@�\=lf�?.            �P@������������������������       �        $             K@�       �                    �?$�q-�?
             *@�       �                    �B@z�G�z�?             @������������������������       �                      @�       �                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       
             �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�       �       
             �?$���}��?`            �c@�       �       	          `ff@θ	j*�?             J@�       �                   0c@nM`����?             G@������������������������       �                     @�       �       	             �?������?            �D@�       �                    �?؇���X�?             <@������������������������       �                     .@�       �                    �?�	j*D�?             *@�       �       	          833�?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   `l@�n_Y�K�?
             *@�       �                   e@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?և���X�?             @������������������������       �                     @�       �                   �]@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       	             @�϶O'3�?A            @Z@�       �                    �?.p����??            @Y@�       �                   Pm@��
ц��?             :@�       �                   pe@d}h���?             ,@������������������������       �                     &@������������������������       �                     @�       �       	          pff�?      �?	             (@�       �                   �c@"pc�
�?             &@������������������������       �                     @�       �                    �?      �?              @�       �                   �c@      �?             @������������������������       �                     �?�       �                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   �l@Х-��ٹ?.            �R@������������������������       �                    �A@�       �                    �?ףp=
�?             D@�       �                    c@"pc�
�?	             &@������������������������       �                      @�       �                   t@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   pn@ 	��p�?             =@�       �                   0n@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     8@������������������������       �                     @�t�b�G     h�h(h+K ��h-��R�(KK�KK��h_�B0       Px@     ��@     �i@     �|@     �J@     �y@     �G@     py@      6@      A@      1@      ,@      *@      �?      *@                      �?      @      *@       @      (@       @      @      �?      @              @      �?              �?                      "@       @      �?              �?       @              @      4@      @      @      @                      @      �?      0@              .@      �?      �?              �?      �?              9@     Pw@      6@      n@      &@     �g@      @      4@      @       @      @       @      @                       @              @              (@      @     `e@      @     �c@             �J@      @     �Z@      @     �P@       @               @     �P@       @      4@       @      @       @      �?              �?       @                      @              .@              G@              D@      @      (@              $@      @       @      @                       @      &@     �H@      &@      ?@      @      @      @              @      @      @      �?       @      �?              �?       @               @                      @      @      9@      �?      5@      �?      @              @      �?                      2@      @      @      �?      @      �?                      @       @                      2@      @     �`@       @      `@      �?      `@             @_@      �?      @              @      �?              �?      �?              �?      �?              �?      @      �?                      @      @      @      @               @      @               @       @       @       @                       @     @c@     �G@     �a@      9@     �F@      3@      @      *@       @              @      *@      @      @      @       @       @       @       @                       @       @              �?      @              @      �?                       @      C@      @     �B@      @      ?@              @      @      @      @      @                      @      @              �?      @      �?                      @     �W@      @      ;@      @      6@              @      @      @       @      @              �?       @               @      �?                      @      Q@              ,@      6@      @      �?              �?      @              @      5@      @      *@      @      @      @       @      @              @       @               @      @                       @              "@               @     �f@     �Q@     �T@      ,@      @      @      @      �?      @              �?      �?      �?                      �?      �?      @              @      �?      �?              �?      �?              S@      "@      R@      @      @      @      @      �?      @                      �?      �?       @      �?                       @     �P@      �?      K@              (@      �?      @      �?       @               @      �?              �?       @               @              @      @      @                      @      Y@     �L@      1@     �A@      1@      =@      @              (@      =@      @      8@              .@      @      "@      @      @      @                      @              @       @      @      @      �?      @                      �?      @      @              @      @      �?              �?      @                      @     �T@      6@     �T@      2@      (@      ,@      @      &@              &@      @              "@      @      "@       @      @              @       @       @       @              �?       @      �?       @                      �?      @                      �?     �Q@      @     �A@              B@      @      "@       @       @              �?       @               @      �?              ;@       @      @       @      @                       @      8@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�@ehG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM	hwh(h+K ��h-��R�(KM	��h~�B�9         �                    �?(@n��?J           ��@       y                    �?>��C��?:           �}@       N       
             �?��.�"*�?�            u@       !                    �?6YE�t�?�            �l@                          `p@�k��(A�?*            �M@                           @L@x�����?            �C@������������������������       �                     1@       	                    �?���|���?             6@������������������������       �                      @
                          P`@և���X�?
             ,@                           �Q@      �?              @                          �_@؇���X�?             @������������������������       �                     @                           �P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @                          �`@�G�z��?             4@                           �?�n_Y�K�?	             *@                            Q@�<ݚ�?             "@                          �c@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?                          �e@      �?             @������������������������       �                     @������������������������       �                     �?                           �J@؇���X�?             @������������������������       �                     @               	          033@      �?             @������������������������       �                     �?������������������������       �                     @"       K                   �u@���W���?v            �e@#       2                    �? rc����?r            `d@$       %                   @[@X�Cc�?             ,@������������������������       �                      @&       1                   �a@�q�q�?             (@'       (                   �g@X�<ݚ�?             "@������������������������       �                     �?)       0                   �`@      �?              @*       -                    �?�q�q�?             @+       ,                   �^@      �?             @������������������������       �                     �?������������������������       �                     @.       /                    `@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @3       4                   �U@p���?f            �b@������������������������       �                      @5       B                   Xp@@9G��?e            `b@6       7                   pa@`Ql�R�?C            �W@������������������������       �        %            �G@8       A       	             �?`�q�0ܴ?            �G@9       >                   �a@���}<S�?             7@:       =                    �L@r�q��?             @;       <                     J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @?       @                    �D@�IєX�?             1@������������������������       �                     �?������������������������       �                     0@������������������������       �                     8@C       H                   �b@�NW���?"            �J@D       G                   �Z@ �q�q�?              H@E       F       	          433�?      �?	             0@������������������������       �                      @������������������������       �                     ,@������������������������       �                     @@I       J                    �?���Q��?             @������������������������       �                      @������������������������       �                     @L       M                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @O       x                   �u@H(���o�?D            �Z@P       _                   �b@X&$�E�?@            �X@Q       V       	          ����?����X�?%             L@R       S                    �?Pa�	�?            �@@������������������������       �                     ?@T       U                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?W       ^                    c@�LQ�1	�?             7@X       ]                    �?����X�?             5@Y       Z                   @[@���Q��?             $@������������������������       �                     @[       \       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                      @`       s                   Hq@X��ʑ��?            �E@a       b                    �?     ��?             @@������������������������       �                      @c       f                    �?r�q��?             8@d       e                    ]@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @g       p                   �l@��S���?
             .@h       i                    �G@�q�q�?             "@������������������������       �                     @j       k                   `@���Q��?             @������������������������       �                      @l       m                    �M@�q�q�?             @������������������������       �                     �?n       o                   `Y@      �?              @������������������������       �                     �?������������������������       �                     �?q       r                    �J@r�q��?             @������������������������       �                     @������������������������       �                     �?t       u                   �r@"pc�
�?             &@������������������������       �                     @v       w                   (t@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @z       �                   �v@�wY;��?V             a@{       �       
             �?�t:ɨ�?R            �`@|       }                     R@���1��?A            �Z@������������������������       �        ?             Z@~                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @[@�J�4�?             9@������������������������       �        
             .@�       �       	          433�?���Q��?             $@�       �                    �H@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �\@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �|@      �?             @������������������������       �                      @������������������������       �                      @�       �       
             �?�ωf�?           �{@�       �                    �?П[;U��?f            �e@�       �                   �Q@4�E��
�?>             Z@�       �       
             �?���y4F�?             3@������������������������       �                     �?�       �                   �c@r�q��?
             2@�       �                    @      �?	             0@�       �                    �K@ףp=
�?             $@������������������������       �                     @�       �                   `X@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �n@�ĚpF�?3            @U@�       �                    �?��6}��?$            �N@�       �       	          ���@��k=.��?            �G@�       �                    �?���V��?            �F@������������������������       �                     4@�       �                    �? �o_��?             9@�       �       	          hff�?�8��8��?             (@������������������������       �                     $@�       �                     G@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �\@��
ц��?
             *@������������������������       �                      @�       �       	            �?���|���?	             &@�       �                    �?      �?             @�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     @�       �                   0j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   @l@      �?             ,@�       �                    �K@      �?              @������������������������       �                      @������������������������       �                     @�       �       	          ����?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �p@      �?             8@������������������������       �                     @�       �       	          ����?�q�q�?             2@�       �                   hq@����X�?             @������������������������       �                     �?�       �                   �s@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   `c@�C��2(�?             &@������������������������       �                     @�       �                    �?r�q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?���L��?(            �Q@�       �                   �\@���!pc�?             &@������������������������       �                     @�       �       
             �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   @Z@@�r-��?!            �M@������������������������       �                     �?�       �                    �D@\-��p�?              M@������������������������       �                     @�       �                    �N@�C��2(�?            �K@�       �                    @N@��hJ,�?             A@�       �                   @e@@4և���?             <@�       �                    �?`2U0*��?             9@�       �       	             �?�C��2(�?             &@������������������������       �                     @�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             ,@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �        
             5@�                           �?$�T@	��?�            �p@�       �                    �?�&/�E�?�             o@�       �                    �?@�0�!��?             A@������������������������       �                     "@�       �                   �c@�+e�X�?             9@�       �                   �k@��2(&�?             6@������������������������       �                     $@�       �                     L@      �?             (@������������������������       �                      @�       �                     P@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	            �?PԱ�l�?�            �j@������������������������       �        q             f@�       �                   pa@���y4F�?             C@������������������������       �                     .@�       �                    �I@�LQ�1	�?             7@������������������������       �                     @�       �       	          033�?      �?
             0@�       �                    @�z�G��?             $@�       �                   b@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    U@r�q��?             @������������������������       �                     �?������������������������       �                     @            	          ����?�û��|�?             7@                        �X@@�0�!��?             1@������������������������       �                     �?                         �?      �?             0@                         �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     $@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM	KK��h_�B�       @{@      ~@     �[@     �v@     �Y@     @m@     �A@     �h@      1@      E@       @      ?@              1@       @      ,@               @       @      @       @      @      �?      @              @      �?       @      �?                       @      �?              @              "@      &@       @      @      @       @      @      �?      @                      �?              �?      �?      @              @      �?              �?      @              @      �?      @      �?                      @      2@     @c@      *@     �b@      @      "@               @      @      @      @      @      �?              @      @       @      @      �?      @      �?                      @      �?      �?              �?      �?               @                      @       @     �a@       @              @     �a@       @      W@             �G@       @     �F@       @      5@      �?      @      �?       @               @      �?                      @      �?      0@      �?                      0@              8@      @     �H@       @      G@       @      ,@       @                      ,@              @@       @      @       @                      @      @      @              @      @              Q@      C@     �N@      C@      D@      0@      @@      �?      ?@              �?      �?              �?      �?               @      .@      @      .@      @      @              @      @      �?      @                      �?              &@       @              5@      6@      3@      *@       @              &@      *@      @      @              @      @              @       @      @      @      @               @      @               @       @      �?      �?              �?      �?      �?                      �?      �?      @              @      �?               @      "@              @       @       @       @                       @      @              @      `@      @     �_@      �?     �Z@              Z@      �?       @      �?                       @      @      5@              .@      @      @      @       @               @      @              �?      @      �?                      @       @       @       @                       @     `t@     �]@     �S@      X@     �N@     �E@      @      .@      �?              @      .@      �?      .@      �?      "@              @      �?      @      �?                      @              @       @             �L@      <@     �F@      0@      C@      "@      C@      @      4@              2@      @      &@      �?      $@              �?      �?      �?                      �?      @      @               @      @      @      �?      @      �?      �?              �?      �?                       @      @      �?      @              �?      �?              �?      �?                       @      @      @       @      @       @                      @      @      �?              �?      @              (@      (@              @      (@      @       @      @      �?              �?      @              @      �?              $@      �?      @              @      �?       @      �?              �?       @              @              1@     �J@       @      @      @              �?      @      �?                      @      "@      I@      �?               @      I@      @              @      I@      @      =@       @      :@      �?      8@      �?      $@              @      �?      @      �?                      @              ,@      �?       @               @      �?              @      @              @      @                      5@      o@      7@     @m@      ,@      <@      @      "@              3@      @      3@      @      $@              "@      @       @              �?      @              @      �?                      @     �i@       @      f@              >@       @      .@              .@       @      @               @       @      @      @      @       @               @      @                      @      @      �?              �?      @              ,@      "@      ,@      @              �?      ,@       @      @       @               @      @              $@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��2hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK酔h~�B�2         X                   �`@��e�B��?>           ��@       '       	             �?�������?           �x@              
             �?���-��?`            `b@                            F@ 7���B�?3            @T@                          �`@      �?             @������������������������       �                     @������������������������       �                     �?              
             �?�g<a�?/            @S@	       
                    \@      �?              @������������������������       �                     �?������������������������       �                     �?                           `@�}��L�?-            �R@                           �O@Pa�	�?            �@@������������������������       �                     =@                          �X@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     E@                          `T@6YE�t�?-            �P@                           �?և���X�?             ,@                           @M@�q�q�?	             "@              	          @33�?      �?             @������������������������       �                      @������������������������       �                      @              	          ����?z�G�z�?             @              	             п      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @       $                    @P@ ��WV�?"             J@        !                   `c@@�E�x�?            �H@������������������������       �                    �E@"       #                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @%       &                     Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @(       K                   @r@��仞�?�             o@)       .                    �?b �57�?�            �i@*       -                     P@և���X�?             ,@+       ,       	          ����?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @/       H                    �Q@ �q�q�?}             h@0       C       
             �?(��m,��?w            @g@1       8                    @O@�h����?l             e@2       3                   `b@���б�?T            �`@������������������������       �        ?             Y@4       5                    �?��?^�k�?            �A@������������������������       �                      @6       7                     F@ 7���B�?             ;@������������������������       �                     �?������������������������       �                     :@9       >                    �O@�FVQ&�?            �@@:       =       
             �?z�G�z�?             @;       <                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @?       B                   `Y@h�����?             <@@       A                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     :@D       E                    _@�<ݚ�?             2@������������������������       �                     &@F       G                    �?և���X�?             @������������������������       �                     @������������������������       �                     @I       J                   `c@r�q��?             @������������������������       �                     @������������������������       �                     �?L       Q                    �?&^�)b�?            �E@M       P                   �t@�q�q�?             (@N       O                    �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @R       W       	             �?�g�y��?             ?@S       T                    �K@�����H�?             "@������������������������       �                     @U       V                   xs@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     6@Y       �                    �?o����?8           P�@Z       �       	          ����?H��%�R�?u            �h@[       \                   @E@I� ��?9             W@������������������������       �                     *@]       �                    �?�;u�,a�?2            �S@^       {       	          ����?b����?(            �O@_       f                    �?(옄��?             G@`       e                   pf@և���X�?             @a       d                    �?�q�q�?             @b       c                    �K@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     �?g       z                    �?��Zy�?            �C@h       y                    �?D�n�3�?             C@i       j                   �g@��J�fj�?            �B@������������������������       �                     @k       l                   0a@�'�=z��?            �@@������������������������       �                      @m       n       
             �?`՟�G��?             ?@������������������������       �                     $@o       p                   �i@��s����?             5@������������������������       �                      @q       x                   @b@�KM�]�?             3@r       s                    �?�X�<ݺ?             2@������������������������       �                     @t       w                    ]@��S�ۿ?	             .@u       v                    �G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?|       �       
             �?�IєX�?
             1@}       ~                   �^@؇���X�?             @������������������������       �                     @       �                   pd@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                     F@      �?
             0@������������������������       �                     @�       �                    b@�q�q�?             (@�       �                    �?�����H�?             "@�       �                   �n@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       
             �?��s�n�?<             Z@�       �                   `b@X��%�?/            �U@�       �                   �a@XB���?             M@�       �                    �? >�֕�?            �A@�       �                    \@$�q-�?             :@�       �                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     7@������������������������       �                     "@������������������������       �                     7@�       �                   �Z@ܷ��?��?             =@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?�>����?             ;@������������������������       �                     $@�       �       	          ����?�t����?
             1@������������������������       �                     �?�       �                   Pc@      �?	             0@�       �                    �?r�q��?             @�       �                   p@�q�q�?             @������������������������       �                     �?�       �                    c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     1@�       �                   �O@8��P�?�            `t@�       �       	             �?X�Cc�?	             ,@�       �                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          033@�Rez��?�            �s@�       �       
             �?��NX��?�            �r@�       �                    �?�q�q�?0            �S@�       �                   �_@���BK�?*            �Q@�       �                   �d@l��\��?             A@�       �                   @q@`Jj��?             ?@�       �       	          ����?h�����?             <@������������������������       �                     3@�       �                    �?�����H�?             "@������������������������       �                     @�       �                   `b@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   `k@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @P@��J�fj�?            �B@�       �                    `@���|���?            �@@������������������������       �                      @�       �                   �o@�4�����?             ?@�       �                    �B@"pc�
�?             6@������������������������       �                     �?�       �                    �H@؇���X�?             5@������������������������       �                      @�       �                   @f@�θ�?
             *@������������������������       �                     �?�       �                    �I@r�q��?	             (@������������������������       �                     �?�       �       	          ����?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �       	          ����?�q�q�?             "@������������������������       �                     @�       �                     @      �?             @������������������������       �                      @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       	            �?����>4�?�             l@������������������������       �        k            �f@�       �                    �?��Y��]�?            �D@�       �                   �_@г�wY;�?             A@�       �                   �^@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?������������������������       �                     5@������������������������       �                     @�       �                   g@�z�G��?             $@�       �                    �?      �?              @�       �       
             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@     @T@     �s@     �M@      V@      @     �S@      �?      @              @      �?               @     �R@      �?      �?              �?      �?              �?     �R@      �?      @@              =@      �?      @              @      �?                      E@      L@      $@      @       @      @      @       @       @       @                       @      @      �?      �?      �?      �?                      �?      @                      @      I@       @      H@      �?     �E@              @      �?              �?      @               @      �?              �?       @              6@     `l@      ,@      h@      @       @       @       @       @                       @      @               @      g@      @     `f@      @     �d@      �?     �`@              Y@      �?      A@               @      �?      :@      �?                      :@       @      ?@      �?      @      �?      �?              �?      �?                      @      �?      ;@      �?      �?      �?                      �?              :@      @      ,@              &@      @      @              @      @              �?      @              @      �?               @     �A@      @      @      @      �?      @                      �?              @      �?      >@      �?       @              @      �?      @              @      �?                      6@     �t@     �g@      I@     @b@     �F@     �G@              *@     �F@      A@     �D@      6@      9@      5@      @      @       @      @       @       @       @                       @               @      �?              6@      1@      6@      0@      5@      0@      @              1@      0@               @      1@      ,@              $@      1@      @               @      1@       @      1@      �?      @              ,@      �?      �?      �?      �?                      �?      *@                      �?      �?                      �?      0@      �?      @      �?      @              @      �?      @                      �?      $@              @      (@              @      @       @      �?       @      �?       @      �?                       @              @      @              @     �X@      @     �T@       @      L@       @     �@@       @      8@       @      �?       @                      �?              7@              "@              7@      @      :@      �?      �?      �?                      �?       @      9@              $@       @      .@      �?              �?      .@      �?      @      �?       @              �?      �?      �?              �?      �?                      @              $@              1@     �q@     �E@      @      "@      @      @              @      @                      @     `q@      A@     0q@      ;@      J@      :@      J@      3@      ?@      @      =@       @      ;@      �?      3@               @      �?      @               @      �?       @                      �?       @      �?              �?       @               @      �?       @                      �?      5@      0@      5@      (@               @      5@      $@      2@      @              �?      2@      @       @              $@      @              �?      $@       @              �?      $@      �?              �?      $@              @      @              @      @      �?       @              �?      �?              �?      �?                      @              @     �k@      �?     �f@              D@      �?     �@@      �?      (@      �?      (@                      �?      5@              @              @      @      �?      @      �?      @      �?                      @              @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ(��uhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�Bx6         �                    �?~jÚʞ�?2           ��@       �                   �f@λ�@��?2            @       6       	          ����?���^��?-           P~@       +                    �?���ѽ��?f             d@       "                    �?.T�߸��?P             _@       	                   @E@Ї?��f�?7            @U@                            G@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@
              
             �?���o,��?0            @R@              	          ����?"pc�
�?             6@������������������������       �                     2@������������������������       �                     @                          @b@�:�]��?!            �I@                          �l@`�q�0ܴ?            �G@������������������������       �                     9@                           �?�C��2(�?             6@������������������������       �                     $@                          @Z@r�q��?	             (@������������������������       �                     �?                          @^@�C��2(�?             &@                           �?z�G�z�?             @                          �[@      �?             @������������������������       �                      @                           @G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �E@      �?             @������������������������       �                     �?        !                    e@�q�q�?             @������������������������       �                     �?������������������������       �                      @#       $                    a@�ݜ�?            �C@������������������������       �                     2@%       (                   �b@���N8�?             5@&       '       
             �?r�q��?             2@������������������������       �                     .@������������������������       �                     @)       *                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?,       1                    �?�L���?            �B@-       .                   0a@(;L]n�?             >@������������������������       �                     9@/       0                   @a@z�G�z�?             @������������������������       �                     @������������������������       �                     �?2       3       
             �?����X�?             @������������������������       �                     @4       5                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?7       R                    �?М-�:�?�            @t@8       K                   xr@\-��p�?0            �U@9       H                   Pe@��S�ۿ?*            �R@:       G                    �?F��}��?(            @R@;       F                   c@��� ��?             ?@<       =                   �U@ףp=
�?             >@������������������������       �                     �?>       E       	          ����? 	��p�?             =@?       @                    �?r�q��?             (@������������������������       �                     �?A       B       	          ����?�C��2(�?             &@������������������������       �                     "@C       D                    @G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     1@������������������������       �                     �?������������������������       �                     E@I       J                    �?      �?              @������������������������       �                     �?������������������������       �                     �?L       O                    �?�q�q�?             (@M       N                   y@r�q��?             @������������������������       �                     @������������������������       �                     �?P       Q       	          @33�?�q�q�?             @������������������������       �                      @������������������������       �                     @S       ~       
             �?@Ix�<��?�            �m@T       }                    �?���O�?�            `k@U       |                    �N@ 	��p�?b             b@V       W                   e@4և����?N             \@������������������������       �                     4@X       q       	          ����?�q��/��?B             W@Y       Z                   �g@      �?             @@������������������������       �                      @[       p                   �e@z�G�z�?             >@\       ]       
             �?д>��C�?             =@������������������������       �                     @^       _       	          ����?��<b���?             7@������������������������       �                     �?`       a                    �G@"pc�
�?             6@������������������������       �                     @b       g                   �l@���y4F�?             3@c       f                    `@���Q��?             @d       e                   �_@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?h       o                    _@؇���X�?             ,@i       j                   @_@����X�?             @������������������������       �                     �?k       n                   �r@r�q��?             @l       m                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?r       w       	          033@(;L]n�?(             N@s       v       	          ���@����?�?            �F@t       u                    c@�g�y��?             ?@������������������������       �                     >@������������������������       �                     �?������������������������       �                     ,@x       {                    �J@��S�ۿ?             .@y       z                    @J@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                    �@@������������������������       �        (            �R@       �       	             �?r�q��?             2@�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �^@��S�ۿ?             .@�       �       	             �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?��^�_�?            `z@�       �       
             �?8�C�M�?�            �q@�       �                    �?��Q:��?&            �M@�       �                    �K@     ��?             0@�       �                    �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                    `P@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?�%^�?            �E@�       �                   xq@�z�G��?             $@������������������������       �                     @������������������������       �                     @�       �                     E@<���D�?            �@@�       �                    �C@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �^@��a�n`�?             ?@�       �                    �?      �?	             (@�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �Z@z�G�z�?             $@�       �                    V@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �        
             3@�       �                   �s@P�Lt�<�?�            �l@�       �                   c@�O4R���?{            �j@�       �                     R@�94�s0�?B            �\@�       �                    �G@P�Lt�<�?A            �\@�       �                    �?@4և���?             E@������������������������       �                     9@�       �                   �b@@�0�!��?	             1@������������������������       �                     ,@������������������������       �                     @������������������������       �        ,             R@������������������������       �                     �?������������������������       �        9            @X@�       �                   �c@      �?
             0@�       �                    `@      �?              @������������������������       �                     @�       �                   0c@      �?             @������������������������       �                     �?�       �                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �b@|��?���?U            �`@�       �                    �?�q�q�?1             R@�       �                     I@<|ۤ$�?%            �K@�       �                    �?8�Z$���?	             *@������������������������       �                     �?�       �                   0b@�8��8��?             (@������������������������       �                     $@�       �       	          `ff@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?             E@������������������������       �                      @�       �                   �e@h+�v:�?             A@�       �       
             �?�c�Α�?             =@�       �                   �r@���B���?             :@�       �                    b@      �?             8@�       �                    @K@@�0�!��?             1@������������������������       �                      @�       �                   �b@��S�ۿ?	             .@������������������������       �                     (@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �a@�IєX�?             1@������������������������       �        	             ,@�       �       	          033�?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �q@�b��-8�?$            �O@�       �       	             @�q�q�?            �I@�       �       	          pff�?>A�F<�?             C@�       �                    �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �O@؇���X�?            �A@�       �       	          ����?�t����?             A@�       �                     M@�>����?             ;@�       �                    �? �q�q�?             8@�       �       	          033�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     5@�       �                    a@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @H@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �B@�θ�?             *@�       �                   �e@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     (@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@     �W@     y@     @U@      y@      N@     @Y@     �L@     �P@      J@     �@@      �?      &@      �?                      &@     �I@      6@      @      2@              2@      @             �G@      @     �F@       @      9@              4@       @      $@              $@       @              �?      $@      �?      @      �?      @      �?       @              �?      �?      �?                      �?      �?              @               @       @              �?       @      �?              �?       @              @      A@              2@      @      0@      @      .@              .@      @               @      �?       @                      �?      @      A@      �?      =@              9@      �?      @              @      �?               @      @              @       @      �?       @                      �?      9@     �r@      (@     �R@      @     �Q@      @     @Q@      @      ;@      @      ;@      �?               @      ;@       @      $@      �?              �?      $@              "@      �?      �?              �?      �?                      1@      �?                      E@      �?      �?      �?                      �?      @      @      @      �?      @                      �?       @      @       @                      @      *@      l@      $@      j@      $@     �`@      $@     �Y@              4@      $@     �T@       @      8@       @              @      8@      @      8@              @      @      2@      �?              @      2@              @      @      .@       @      @      �?      @      �?                      @      �?               @      (@       @      @      �?              �?      @      �?       @               @      �?                      @              @      �?               @      M@      �?      F@      �?      >@              >@      �?                      ,@      �?      ,@      �?      @              @      �?                      "@             �@@             �R@      @      .@       @      �?              �?       @              �?      ,@      �?      @              @      �?                      "@      $@      �?      @              @      �?      @                      �?     �s@      [@     �n@     �E@      6@     �B@      &@      @      "@      �?      "@                      �?       @      @              @       @              &@      @@      @      @      @                      @      @      =@      �?      �?              �?      �?              @      <@      @      "@      �?      �?      �?                      �?       @       @       @      �?              �?       @                      @              3@     �k@      @      j@      @     �[@      @     �[@      @     �C@      @      9@              ,@      @      ,@                      @      R@                      �?     @X@              ,@       @      @       @      @               @       @              �?       @      �?              �?       @               @             �Q@     @P@      8@      H@      7@      @@       @      &@      �?              �?      &@              $@      �?      �?      �?                      �?      5@      5@       @              *@      5@       @      5@      @      5@      @      5@      @      ,@       @              �?      ,@              (@      �?       @      �?                       @              @       @              @              @              �?      0@              ,@      �?       @               @      �?              G@      1@      A@      1@      ?@      @      �?       @      �?                       @      >@      @      >@      @      9@       @      7@      �?       @      �?              �?       @              5@               @      �?              �?       @              @       @               @      @                      �?      @      $@      @       @               @      @                       @      (@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�ChG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKh~�BH4         �                    �?Ly�'^��?2           ��@       Y       
             �?ƆQ����?*           �~@       R                   �u@�KM�]�?�            `u@       	                    b@������?�            �t@                           @O@���E�?7            �U@������������������������       �        +            @Q@              
             �?�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@
                          @Z@�L�� ��?�            �n@                           �B@      �?             @������������������������       �                     �?������������������������       �                     @       #                    �?���(\��?�             n@                          �g@�	j*D�?            �C@������������������������       �                     @                           �J@4�2%ޑ�?            �A@                          @[@�q�q�?             "@������������������������       �                      @                           @I@؇���X�?             @������������������������       �                     @                          �q@      �?              @������������������������       �                     �?������������������������       �                     �?       "                   �`@$�q-�?             :@       !                   �`@"pc�
�?             &@                           @L@      �?             @������������������������       �                     �?                           �?�q�q�?             @������������������������       �                     �?               	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     .@$       Q                   �e@t�e�í�?u             i@%       D                   Pb@�-m7"C�?t            �h@&       '                    �?�f"Nf�?h             f@������������������������       �                     D@(       -                   @X@A_�&�?Q             a@)       *                    @K@�<ݚ�?             "@������������������������       �                     @+       ,                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @.       1                   pe@     �?L             `@/       0                    _@�q�q�?             @������������������������       �                     @������������������������       �                      @2       3                   0p@�]0��<�?H            �^@������������������������       �        *            �O@4       C                    �R@ ,��-�?            �M@5       <                   �p@�8���?             M@6       7       	          ����?      �?              @������������������������       �                      @8       9       	          ����?�q�q�?             @������������������������       �                     �?:       ;                     M@z�G�z�?             @������������������������       �                     �?������������������������       �                     @=       B                    �?p���?             I@>       A                   @_@      �?             @@?       @       	             �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     8@������������������������       �                     2@������������������������       �                     �?E       P                   pb@�GN�z�?             6@F       G                   �h@     ��?
             0@������������������������       �                      @H       K                   Pq@d}h���?	             ,@I       J       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @L       M                   �b@�����H�?             "@������������������������       �                     @N       O                    �O@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @S       T                     L@�eP*L��?             &@������������������������       �                     @U       V                   `v@r�q��?             @������������������������       �                     @W       X                    @O@�q�q�?             @������������������������       �                      @������������������������       �                     �?Z       �                   0f@��-*��?W            @b@[       �                    �?���nU��?P            ``@\       q                   pc@���@M^�?;            @W@]       f                    �?      �?&             N@^       _       	          ����?$G$n��?            �B@������������������������       �                     8@`       c                   �m@�n_Y�K�?             *@a       b                   ``@      �?              @������������������������       �                      @������������������������       �                     @d       e                    �?���Q��?             @������������������������       �                     @������������������������       �                      @g       h                   �[@\X��t�?             7@������������������������       �                     @i       j                   �]@�����?             3@������������������������       �                     @k       l       	             �?      �?             (@������������������������       �                      @m       p                   �`@���Q��?             $@n       o                   c@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @r       {                    �?���|���?            �@@s       t                   �i@�eP*L��?             6@������������������������       �                     @u       v                    �G@X�<ݚ�?             2@������������������������       �                      @w       z                    �L@z�G�z�?             $@x       y                    m@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @|       }                   �^@"pc�
�?             &@������������������������       �                     �?~                           @K@ףp=
�?             $@������������������������       �                     @�       �                    h@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   ``@�KM�]�?             C@������������������������       �                     =@�       �                   �a@X�<ݚ�?             "@�       �                   @[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     .@�       �       
             �?�8�0�|�?           �z@�       �                   �b@W����?[             b@�       �                    �?�8=�?B            �Y@�       �                    @N@d}h���?             ,@������������������������       �                     $@�       �                    �?      �?             @�       �                    @Q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?ą%�E�?:            @V@�       �                   �l@�q�q�?             (@�       �                    �?և���X�?             @�       �                    W@z�G�z�?             @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   @Y@XI�~�?/            @S@������������������������       �                      @�       �       
             �?`2U0*��?.            �R@�       �                    d@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                   �[@����e��?(            �P@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        $             N@�       �                    @�ՙ/�?             E@�       �                    �?4�B��?            �B@�       �       	          ����?�������?             A@�       �       	          ����?R���Q�?	             4@�       �                    e@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     (@�       �       	          033�?և���X�?	             ,@�       �                   �q@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?      �?              @�       �                    @L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �G@z�G�z�?             @������������������������       �                     @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @��S�ۿ?�            �q@�       �                    �O@�Xyd�B�?�            �p@�       �                    @L@������?�            �o@�       �                   pf@`׀�:M�?�            �k@�       �                   @[@ 3S6ɓ?w            �i@�       �                   �Z@�FVQ&�?
            �@@������������������������       �                     9@�       �                   �o@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �        m            �e@�       �                    �?�IєX�?             1@������������������������       �        	             .@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �L@�r����?             >@�       �       	          pff�?և���X�?             @�       �                   Hp@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�nkK�?             7@�       �                    �?r�q��?             @������������������������       �                      @�       �                   �p@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     1@�       �                     P@j���� �?             1@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �       	          `ff�?      �?	             (@�       �                    �?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                      @�       �                   `Q@     ��?             0@������������������������       �                      @�       �                   Pp@d}h���?             ,@�       �                   �`@8�Z$���?
             *@�       �                    �J@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�t�b�W     h�h(h+K ��h-��R�(KK�KK��h_�B�       �z@     �~@      \@     �w@      B@      s@      ?@     �r@      �?     �U@             @Q@      �?      1@      �?                      1@      >@     �j@      @      �?              �?      @              ;@     �j@      (@      ;@      @               @      ;@      @      @               @      @      �?      @              �?      �?      �?                      �?       @      8@       @      "@       @       @              �?       @      �?      �?              �?      �?      �?                      �?              @              .@      .@     @g@      *@     @g@       @      e@              D@       @      `@       @      @              @       @      �?              �?       @              @     �^@       @      @              @       @              @     �]@             �O@      @     �K@      @     �K@       @      @               @       @      @      �?              �?      @      �?                      @      �?     �H@      �?      ?@      �?      @      �?                      @              8@              2@      �?              @      1@      @      &@       @              @      &@       @      @              @       @              �?       @              @      �?      @              @      �?                      @       @              @      @              @      @      �?      @               @      �?       @                      �?      S@     �Q@     �N@     �Q@     �L@      B@     �F@      .@      @@      @      8@               @      @      @       @               @      @               @      @              @       @              *@      $@              @      *@      @      @              @      @       @              @      @      @       @      @                       @              @      (@      5@      $@      (@              @      $@       @       @               @       @       @      @              @       @                      @       @      "@      �?              �?      "@              @      �?      @              @      �?              @      A@              =@      @      @      @      �?              �?      @                      @      .@             �s@     �]@      G@     �X@      4@     �T@      &@      @      $@              �?      @      �?      �?              �?      �?                       @      "@      T@      @       @      @      @      @      �?      �?      �?      �?                      �?      @                       @              @      @      R@       @              @      R@       @      @              @       @              �?     @P@      �?      @              @      �?                      N@      :@      0@      9@      (@      9@      "@      1@      @      @      @      @                      @      (@               @      @       @      @              @       @              @       @      �?       @      �?                       @      @                      @      �?      @              @      �?      �?      �?                      �?     �p@      3@     �o@      ,@     �n@      @     `k@      @     `i@       @      ?@       @      9@              @       @               @      @             �e@              0@      �?      .@              �?      �?      �?                      �?      :@      @      @      @      �?      @      �?                      @      @              6@      �?      @      �?       @              @      �?      @                      �?      1@              $@      @      �?      @      �?                      @      "@      @      "@      �?      "@                      �?               @      &@      @               @      &@      @      &@       @      @       @      @                       @       @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��?hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B6         �       
             �?�LT ���?B           ��@       a                    �?L�zF�?M           �@                          �f@����X�?�            @j@                           �?�F��O�?+            @R@������������������������       �                    �G@       	       
             �?�θ�?             :@                            P@�q�q�?             @������������������������       �                      @������������������������       �                     �?
                           �?�㙢�c�?             7@              	          ����?      �?             @������������������������       �                      @������������������������       �                      @                           @G@�KM�]�?
             3@                           _@�q�q�?             @������������������������       �                     �?������������������������       �                      @                          �X@      �?             0@                           X@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@       &       	          ����?(����?\             a@                           �?>A�F<�?             C@������������������������       �                     5@                           �?j���� �?             1@                           �?����X�?             @������������������������       �                     �?                          �\@r�q��?             @������������������������       �                     �?������������������������       �                     @        !                    �?z�G�z�?	             $@������������������������       �                     �?"       #                   @b@�����H�?             "@������������������������       �                     @$       %                   0c@      �?             @������������������������       �                     �?������������������������       �                     @'       H                    �?>����?@            �X@(       -                   @^@���h%��?+            �O@)       *                    �?ףp=
�?             4@������������������������       �        	             .@+       ,                   8w@���Q��?             @������������������������       �                     @������������������������       �                      @.       G                   �a@�K��&�?            �E@/       4                   �\@     ��?             @@0       1                   p@      �?              @������������������������       �                     @2       3                   8r@      �?             @������������������������       �                      @������������������������       �                      @5       6                   �k@�q�q�?             8@������������������������       �                      @7       >                    �?      �?             0@8       9       	          ����?�q�q�?	             "@������������������������       �                      @:       =       	          ����?؇���X�?             @;       <                   xu@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @?       F                   �_@����X�?             @@       E                   pc@���Q��?             @A       D                    �?�q�q�?             @B       C                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     &@I       R                   �b@      �?             B@J       Q                    @$�q-�?             *@K       L                    �?r�q��?             @������������������������       �                      @M       P                    @Q@      �?             @N       O                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @S       X                   �l@�LQ�1	�?             7@T       U                    b@�C��2(�?             &@������������������������       �                     @V       W                    @      �?             @������������������������       �                     �?������������������������       �                     @Y       Z                   �m@�q�q�?             (@������������������������       �                     @[       `       	          ���@����X�?             @\       ]                   �d@      �?             @������������������������       �                     �?^       _       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @b       c                   �U@���Lͩ�?�            �r@������������������������       �                      @d       �                   �b@�
�@c�?�            �r@e       �                    �?dkRk?�?�            pq@f       �       	          ����?�C��2(�?�            �h@g       �                   �s@�ȼB���?N            �[@h       {                    �?      �?G             Z@i       j       	             �?p`q�q��?5            �S@������������������������       �                     3@k       n       	          ����?�?�P�a�?'             N@l       m                   �\@�q�q�?             @������������������������       �                      @������������������������       �                     @o       p                    �?�X�<ݺ?$             K@������������������������       �                     2@q       v       	          033�?�8��8��?             B@r       u                    �? �q�q�?             8@s       t                   �m@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@w       x                   �c@r�q��?             (@������������������������       �                     @y       z                   �_@����X�?             @������������������������       �                     @������������������������       �                      @|       }                   `X@�+e�X�?             9@������������������������       �                      @~                           �H@�㙢�c�?             7@������������������������       �                     �?�       �                   0a@��2(&�?             6@�       �       	          ����?�}�+r��?             3@�       �                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                     "@�       �                    `@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @M@և���X�?             @�       �                   �Y@�q�q�?             @������������������������       �                      @�       �                    �?      �?             @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    �J@�d���??            �U@�       �                    �?�C��2(�?             6@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �k@P���Q�?             4@�       �                   Pb@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             .@������������������������       �        .            @P@�       �                    `P@ �)���?.            @T@������������������������       �        (            �Q@�       �                    ]@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                    �?p�ݯ��?
             3@�       �                    @�q�q�?             (@�       �                    �?���|���?             &@�       �       	             �?      �?              @�       �                   c@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   @E@Қc,���?�            �y@�       �       	            �?��E�B��?            �G@�       �                    �?�q�q�?             2@�       �                    �?և���X�?             ,@�       �                   �b@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     =@�       �       	          033@��h��Q�?�            �v@�       �                    �?LW�S�?�            0v@�       �                    _@����X�?:            �V@�       �                   0q@�X�<ݺ?             B@�       �                   �a@Pa�	�?            �@@������������������������       �        
             3@�       �                    �?@4և���?	             ,@������������������������       �                     @�       �                    �F@�����H�?             "@������������������������       �                     @�       �                    �G@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    t@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   pc@ؓ��M{�?%            �K@�       �                    �?������?             >@������������������������       �                     1@�       �                   �p@�n_Y�K�?	             *@�       �                    b@      �?              @������������������������       �                     @�       �                   �_@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��H�}�?             9@�       �                   d@      �?             @������������������������       �                     �?�       �                   pe@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    `@�q�q�?             5@������������������������       �                     @�       �                   �f@j���� �?	             1@�       �                   �c@����X�?             ,@������������������������       �                     �?�       �                    �?�θ�?             *@�       �       	          @33�?      �?              @�       �                   (r@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �g@�t:ɨ�?�            �p@�       �                    @L@������?�            Pp@������������������������       �        z            �i@�       �                    �M@X�;�^o�?"            �K@�       �                   0b@     ��?             0@�       �                    �?����X�?             @�       �                   �m@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     "@�       �                   `c@�7��?            �C@������������������������       �                     >@�       �                    �?�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp       �y@     �@      V@     `z@      N@     �b@      @     �P@             �G@      @      4@       @      �?       @                      �?      @      3@       @       @               @       @               @      1@      �?       @      �?                       @      �?      .@      �?      @              @      �?                      &@      K@     �T@      @      ?@              5@      @      $@      @       @              �?      @      �?              �?      @               @       @      �?              �?       @              @      �?      @      �?                      @     �G@      J@      4@     �E@       @      2@              .@       @      @              @       @              2@      9@      2@      ,@       @      @              @       @       @       @                       @      0@       @       @               @       @      @      @       @              �?      @      �?       @               @      �?                      @      @       @      @       @      �?       @      �?      �?      �?                      �?              �?       @               @                      &@      ;@      "@      (@      �?      @      �?       @              @      �?       @      �?       @                      �?      �?              @              .@       @      $@      �?      @              @      �?              �?      @              @      @              @      @       @       @       @      �?              �?       @      �?                       @      @              <@      q@       @              :@      q@      3@     @p@      2@     �f@      0@     �W@      *@     �V@      @      R@              3@      @     �J@      @       @               @      @              @     �I@              2@      @     �@@      �?      7@      �?      @      �?                      @              3@       @      $@              @       @      @              @       @              @      3@       @              @      3@      �?              @      3@      �?      2@      �?      "@      �?                      "@              "@       @      �?       @                      �?      @      @       @      @               @       @       @       @      �?       @                      �?              �?      �?               @     @U@       @      4@      �?      �?              �?      �?              �?      3@      �?      @              @      �?                      .@             @P@      �?      T@             �Q@      �?      "@      �?                      "@      @      (@      @      @      @      @      @      @      �?      @      �?                      @      @              @                      �?              @     Pt@     �T@      @     �D@      @      (@      @       @      @      �?      @                      �?              @              @              =@     �s@      E@     �s@      B@     @P@      :@      A@       @      @@      �?      3@              *@      �?      @               @      �?      @              @      �?              �?      @               @      �?              �?       @              ?@      8@      6@       @      1@              @       @      �?      @              @      �?       @               @      �?              @      �?      @                      �?      "@      0@       @       @      �?              �?       @               @      �?              @      ,@              @      @      $@      @      $@      �?              @      $@      @      @      �?      @              @      �?               @                      @      @             �o@      $@     �o@      @     �i@              H@      @      &@      @       @      @      �?      @      �?                      @      �?              "@             �B@       @      >@              @       @      @                       @              @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��hkhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�Bx6         n       	          `ff�?~jÚʞ�?C           ��@       '       
             �?
������?6           @@                          ph@�ZD����?g            @f@                           �?Ћ����?/            �T@                          �Q@      �?              @������������������������       �                     @������������������������       �                      @       	                    @`׀�:M�?*            �R@������������������������       �        (             R@
                           `@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?r�q��?8             X@                           �?4�2%ޑ�?            �A@                           @N@؇���X�?             <@                          `a@�nkK�?
             7@������������������������       �        	             6@������������������������       �                     �?                           �?���Q��?             @������������������������       �                      @������������������������       �                     @                          `c@և���X�?             @������������������������       �                     @������������������������       �                     @       "       	          833�?��6}��?)            �N@       !                    �?Du9iH��?            �E@                             E@ �Cc}�?             <@                           �?      �?              @������������������������       �                     @                          �^@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@������������������������       �                     .@#       $                     J@�E��ӭ�?             2@������������������������       �                     @%       &                    �?�r����?	             .@������������������������       �                     *@������������������������       �                      @(       3                   @E@���!r�?�             t@)       0                    �?և���X�?
             ,@*       /                    �?      �?              @+       ,                   �_@r�q��?             @������������������������       �                     @-       .                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @1       2                    `Q@r�q��?             @������������������������       �                     @������������������������       �                     �?4       g                    �? �Cc}�?�            @s@5       J                    �?��|C_�?�            �q@6       =                    q@l��
I��?"             K@7       <                    _@��hJ,�?             A@8       9                   j@�eP*L��?             &@������������������������       �                     @:       ;                     H@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     7@>       E                   �d@�G�z��?             4@?       D                    v@���!pc�?             &@@       C                   ps@���Q��?             @A       B                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @F       G                   f@�����H�?             "@������������������������       �                     @H       I                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?K       T                    �L@@�?1X�?�            �l@L       S                   `\@���ʄ?~            �h@M       R                    �?      �?             @@N       O                   �k@      �?             @������������������������       �                      @P       Q                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     <@������������������������       �        i            �d@U       b                    @"pc�
�?            �@@V       W                   @Y@�����H�?             ;@������������������������       �                     �?X       Y                    @N@$�q-�?             :@������������������������       �        	             ,@Z       a       	          ����?r�q��?	             (@[       `                   @d@����X�?             @\       _                    �?�q�q�?             @]       ^                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @c       d                   `a@      �?             @������������������������       �                      @e       f                   �k@      �?             @������������������������       �                     @������������������������       �                     �?h       m                    �?���Q��?             9@i       l                   �b@�q�q�?	             .@j       k                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     $@o       �                   Xr@޷��$/�?            z@p       �                    �?��;��?�            �u@q       �                   d@Fx$(�?!             I@r       }                    �?����>�?            �B@s       t                   @X@�>����?             ;@������������������������       �                     �?u       |       	          033�? ��WV�?             :@v       w                    �?ףp=
�?             $@������������������������       �                      @x       {                     L@      �?              @y       z                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     0@~       �       	             �?z�G�z�?	             $@       �                   �`@����X�?             @�       �                   @n@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?�	j*D�?             *@�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �Y@�]ؘw��?�            �r@�       �       	             @����X�?             @�       �                    �G@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   0b@,Ӕ��?�            @r@�       �                    �?`-�I�w�?�            �l@�       �                    �?�?�|�?y             g@�       �                    �?Pa�	�?            �@@������������������������       �                     8@�       �                    `@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       
             �?P�Lt�<�?b             c@�       �       	          ����?`��(�?W            �`@�       �                    �?�>����?             ;@������������������������       �                     3@�       �                    ^@      �?              @������������������������       �                     �?�       �                   �`@؇���X�?             @�       �                   �X@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        C             [@�       �                    c@�t����?             1@������������������������       �                     *@�       �                   �_@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �X@>��C��?            �E@������������������������       �                     @�       �                   pb@z�G�z�?             D@�       �                    @F@�����H�?             B@������������������������       �                      @�       �       
             �?�IєX�?             A@������������������������       �                     >@�       �                    �?      �?             @������������������������       �                     �?�       �                     M@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �       
             �?     ��?'             P@�       �                   `d@RB)��.�?            �E@�       �                   �m@��R[s�?            �A@�       �                   �j@X�<ݚ�?             2@�       �                    �F@"pc�
�?             &@������������������������       �                     �?�       �                    @M@ףp=
�?             $@������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          ���@؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �                    q@�IєX�?
             1@������������������������       �                     $@�       �                    @M@؇���X�?             @������������������������       �                     @�       �                     N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    @D@�G��l��?             5@������������������������       �                     @�       �                   �l@j���� �?
             1@�       �                    @K@�θ�?             *@������������������������       �                      @�       �                   �h@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   c@�q�q�?+            @Q@�       �       
             �?�BbΊ�?#             M@�       �                   @^@4և����?!             L@�       �       	             �?ҳ�wY;�?             A@�       �                   �c@b�2�tk�?             2@�       �                    Z@������?             .@������������������������       �                     @�       �                   �t@���Q��?             $@�       �                    �?      �?              @�       �                   �\@����X�?             @�       �                   �s@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    c@      �?
             0@������������������������       �                     $@�       �       
             �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   �r@���7�?             6@�       �                   ``@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@������������������������       �                      @�       �                    �?���!pc�?             &@�       �                    b@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@     pt@     �e@      G@     �`@      @     �S@       @      @              @       @              �?     @R@              R@      �?      �?      �?                      �?     �E@     �J@      ;@       @      8@      @      6@      �?      6@                      �?       @      @       @                      @      @      @              @      @              0@     �F@      @      D@      @      9@      @      @              @      @      �?              �?      @                      4@              .@      *@      @              @      *@       @      *@                       @     �q@     �D@      @       @      �?      @      �?      @              @      �?      �?      �?                      �?               @      @      �?      @                      �?     0q@     �@@     @p@      7@      C@      0@      =@      @      @      @              @      @      �?              �?      @              7@              "@      &@       @      @       @      @       @      �?       @                      �?               @      @              �?       @              @      �?       @               @      �?             �k@      @     `h@      �?      ?@      �?      @      �?       @              �?      �?      �?                      �?      <@             �d@              ;@      @      8@      @              �?      8@       @      ,@              $@       @      @       @      �?       @      �?      �?      �?                      �?              �?      @              @              @      @       @              �?      @              @      �?              .@      $@      @      $@      @      @              @      @                      @      $@             �T@      u@     �M@      r@      3@      ?@      $@      ;@       @      9@      �?              �?      9@      �?      "@               @      �?      @      �?       @      �?                       @              @              0@       @       @      @       @       @       @       @                       @      @              @              "@      @      �?      @      �?      �?      �?                      �?              @       @              D@     0p@      @       @      @      �?              �?      @                      �?     �A@     p@      .@     �j@      @     �f@      �?      @@              8@      �?       @      �?                       @      @     �b@       @     �`@       @      9@              3@       @      @      �?              �?      @      �?      @      �?                      @              @              [@       @      .@              *@       @       @               @       @              $@     �@@      @              @     �@@      @      @@       @               @      @@              >@       @       @      �?              �?       @      �?                       @      @      �?              �?      @              4@      F@      "@      A@      "@      :@       @      $@       @      "@      �?              �?      "@              @      �?       @               @      �?              @      �?      @                      �?      �?      0@              $@      �?      @              @      �?       @      �?                       @               @      &@      $@      @              @      $@      @      $@               @      @       @      @                       @      @              7@      G@      .@     �E@      *@     �E@      (@      6@      &@      @      &@      @      @              @      @      @       @      @       @      @       @               @      @               @              �?                       @              @      �?      .@              $@      �?      @      �?                      @      �?      5@      �?      �?              �?      �?                      4@       @               @      @       @      �?       @                      �?               @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��6zhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B88         �       	          033�?�m=62}�?J           ��@                          @E@ĳ�&���?7           �~@       
                    �?�*/�8V�?;            �W@       	                    �?��
���?/            �R@                          �Z@�7��?            �C@������������������������       �                     4@                          @\@�KM�]�?             3@������������������������       �                      @������������������������       �                     1@������������������������       �                     B@              
             �?D�n�3�?             3@������������������������       �                     &@������������������������       �                      @       g                    �?�� ��?�             y@       2                    �?�Q�ś�?�            �t@              
             �?��>4և�?:             U@                           �?H�V�e��?             A@                           �?      �?             @������������������������       �                     @������������������������       �                     �?                          �]@�r����?             >@������������������������       �                     @                          �b@�㙢�c�?             7@                           `@�}�+r��?
             3@              	             �?�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     $@                          �k@      �?             @������������������������       �                     �?������������������������       �                     @        +                   �_@H%u��?$             I@!       "                   pl@��<b���?             7@������������������������       �        	             ,@#       *                   �c@X�<ݚ�?             "@$       %                   0m@�q�q�?             @������������������������       �                      @&       '                    �?      �?             @������������������������       �                     �?(       )                    @E@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @,       -                    b@ 7���B�?             ;@������������������������       �                     6@.       /                   �f@z�G�z�?             @������������������������       �                     @0       1                    @J@      �?              @������������������������       �                     �?������������������������       �                     �?3       J       
             �?HP�s��?�            @o@4       E                   `a@���|���?            �@@5       >                   `o@�q�q�?             8@6       =                    @L@�����H�?             2@7       8                    @G@�IєX�?
             1@������������������������       �                     &@9       :                    �?r�q��?             @������������������������       �                     @;       <                     I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �??       @                    �?      �?             @������������������������       �                      @A       B                   �b@      �?             @������������������������       �                      @C       D                   e@      �?              @������������������������       �                     �?������������������������       �                     �?F       I                    �?�<ݚ�?             "@G       H                    �N@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @K       N                    c@�&�� .�?�             k@L       M                   p`@      �?              @������������������������       �                      @������������������������       �                     @O       d                    �? Os���?�             j@P       [                    �?��Μ�V�?w             h@Q       R                   `_@�KM�]�?             3@������������������������       �                     �?S       Z                    �?�X�<ݺ?             2@T       Y                   �d@؇���X�?             @U       V                    @L@�q�q�?             @������������������������       �                     �?W       X                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     &@\       ]                    �?�B:�g�?i            �e@������������������������       �        (             Q@^       _                    �?@䯦s#�?A            �Z@������������������������       �        '            �P@`       c                     H@�(\����?             D@a       b                   @[@���N8�?             5@������������������������       �                     �?������������������������       �                     4@������������������������       �                     3@e       f                   @r@     ��?
             0@������������������������       �        	             *@������������������������       �                     @h       �                   @b@���e��?%            �P@i       v                   ``@z�J��?            �G@j       u                   @d@��+7��?             7@k       r       	          833�?�KM�]�?             3@l       m                     I@�IєX�?             1@������������������������       �                     "@n       o                    �?      �?              @������������������������       �                     @p       q                    �?      �?              @������������������������       �                     �?������������������������       �                     �?s       t                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @w       |                    h@      �?             8@x       y       
             �?����X�?             @������������������������       �                     @z       {                   Pa@      �?             @������������������������       �                      @������������������������       �                      @}       �                   �b@�IєX�?
             1@~                            G@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     *@�       �                    �?�}�+r��?	             3@�       �                     M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@�       �       
             �?r�A�%��?           �z@�       �                    �?J�)m��?�            @w@�       �                    �?����e��?'            �P@�       �                   �`@R�}e�.�?             J@�       �                    �?D�n�3�?             3@�       �                   �`@��S���?	             .@������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?"pc�
�?            �@@�       �                    �?ףp=
�?             >@�       �                    �H@�����H�?             ;@�       �       	             �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�       �                    �?�X�<ݺ?             2@�       �       	          033@�����H�?             "@�       �                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     @������������������������       �                     @�       �                    @؇���X�?	             ,@�       �                   �Z@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@������������������������       �                     @�       �                    �?
����?�             s@�       �                   pr@�������?6            �U@�       �       	          ���@z���=��?1            @S@�       �                   0b@4?,R��?-             R@�       �       	          ����? �q�q�?             H@�       �                    �?���}<S�?             7@�       �                    [@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     *@������������������������       �                     9@�       �                   �`@�q�q�?             8@�       �                    �?��.k���?
             1@�       �       	          033�?�n_Y�K�?             *@������������������������       �                      @�       �                    �?���!pc�?             &@�       �       	          ����?�����H�?             "@������������������������       �                     @�       �                   pd@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �X@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �d@���Q��?             @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   �V@P���Q�?�            �k@������������������������       �                     �?�       �                    _@���O�?�            `k@�       �                    �?�LQ�1	�?"             G@�       �                   �a@�˹�m��?             C@������������������������       �                     >@�       �                    �?      �?              @������������������������       �                      @�       �                    �?r�q��?             @�       �                     D@z�G�z�?             @������������������������       �                     @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �^@      �?              @������������������������       �                     @������������������������       �                     @�       �                   �b@����� �?n            �e@�       �                   �b@ �|ك�?O            �^@������������������������       �        M             ^@�       �                   `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �r@ "��u�?             I@�       �       	          ����?P�Lt�<�?             C@�       �                   �_@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     =@�       �                   �s@r�q��?             (@�       �                   �c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                    �?��B����?%             J@�       �                   �u@�c�Α�?             =@�       �                    �H@�<ݚ�?             ;@�       �                   p`@���Q��?             @�       �                    @F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   �c@��2(&�?             6@�       �                   �^@P���Q�?             4@�       �                   a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@������������������������       �                      @������������������������       �                      @�       �                    �?�㙢�c�?             7@������������������������       �                     "@�       �                    �?����X�?
             ,@�       �                   �e@�����H�?             "@������������������������       �                      @������������������������       �                     �?�                           �M@���Q��?             @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�B       y@     (�@     �s@     @f@      $@      U@       @     @R@       @     �B@              4@       @      1@       @                      1@              B@       @      &@              &@       @              s@     �W@     �q@     �J@     �I@     �@@      @      ;@      @      �?      @                      �?      @      :@              @      @      3@      �?      2@      �?       @               @      �?                      $@      @      �?              �?      @              F@      @      2@      @      ,@              @      @      @       @       @               @       @      �?              �?       @      �?                       @              @      :@      �?      6@              @      �?      @              �?      �?      �?                      �?     �l@      4@      5@      (@      3@      @      0@       @      0@      �?      &@              @      �?      @              �?      �?              �?      �?                      �?      @      @       @              �?      @               @      �?      �?      �?                      �?       @      @       @       @               @       @                      @      j@       @      @       @               @      @             `i@      @     �g@      @      1@       @              �?      1@      �?      @      �?       @      �?      �?              �?      �?              �?      �?              @              &@             �e@      �?      Q@             @Z@      �?     �P@             �C@      �?      4@      �?              �?      4@              3@              *@      @      *@                      @      9@     �D@      8@      7@      @      1@       @      1@      �?      0@              "@      �?      @              @      �?      �?              �?      �?              �?      �?      �?                      �?      @              2@      @       @      @              @       @       @       @                       @      0@      �?      @      �?              �?      @              *@              �?      2@      �?       @      �?                       @              0@     @U@     0u@      M@     �s@      :@      D@      ,@      C@       @      &@       @      @       @                      @              @      @      ;@      @      ;@      @      8@       @      @       @                      @      �?      1@      �?       @      �?      �?      �?                      �?              @              "@              @      @              (@       @      "@       @               @      "@              @              @@      q@      5@     @P@      *@      P@      $@      O@       @      G@       @      5@       @       @       @                       @              *@              9@       @      0@       @      "@      @       @       @              @       @      �?       @              @      �?      @      �?                      @       @              @      �?              �?      @                      @      @       @      �?       @               @      �?               @               @      �?              �?       @              &@      j@      �?              $@      j@      @      D@      @     �A@              >@      @      @       @              �?      @      �?      @              @      �?      �?              �?      �?                      �?      @      @              @      @              @      e@      �?     �^@              ^@      �?       @      �?                       @      @     �G@      �?     �B@      �?       @               @      �?                      =@       @      $@       @       @               @       @                       @      ;@      9@       @      5@      @      5@      @       @      �?       @               @      �?               @              @      3@      �?      3@      �?      �?      �?                      �?              2@       @               @              3@      @      "@              $@      @       @      �?       @                      �?       @      @       @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ|#>~hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�6         �                    �?�~8�e�??           ��@       E       
             �?r�0?��?N           ��@                           �?�K��(��?�            �i@                           �?������?E            �[@              	          ����?�n`���?%             O@                           �?�q�q�?            �@@              	          ����?�q�q�?             "@������������������������       �                      @	       
                   `@؇���X�?             @������������������������       �                     �?������������������������       �                     @                          ``@�q�q�?             8@������������������������       �        	             ,@                          �`@      �?	             $@              	             �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                          �_@XB���?             =@                           �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �        	             3@������������������������       �                     �H@       &                    �?r�q��?>             X@       %                    @8^s]e�?             =@       $                    �?�\��N��?             3@       #                   �e@��.k���?             1@                            �?X�Cc�?	             ,@                          �`@r�q��?             @������������������������       �                     @������������������������       �                     �?!       "                   �b@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     $@'       @                   `a@�#}7��?,            �P@(       1       	          ����?JJ����?            �G@)       *                    �?�z�G��?             4@������������������������       �                     "@+       0                   o@�eP*L��?             &@,       /                   �a@      �?              @-       .                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @2       7                    �?l��
I��?             ;@3       6                    �?���Q��?             @4       5                   @q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @8       ;                    �?�GN�z�?             6@9       :                    �D@      �?	             0@������������������������       �                      @������������������������       �                     ,@<       ?                    `@      �?             @=       >                    _@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @A       D                   @]@P���Q�?             4@B       C                    �R@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             .@F       �                    �?0H�JE)�?�            �t@G       P                   @E@�@z�K9�?�            �q@H       K                    �?ҳ�wY;�?
             1@I       J                   �_@      �?             @������������������������       �                     �?������������������������       �                     @L       M                    �?�n_Y�K�?             *@������������������������       �                     @N       O                    _@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @Q       f                    �?t�e�í�?�            �p@R       a                    @N@8�Z$���?)            @P@S       T                   �c@ܷ��?��?#             M@������������������������       �                    �A@U       Z                    �?��+7��?             7@V       W                    @H@�q�q�?             @������������������������       �                     �?X       Y                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?[       `                   �b@z�G�z�?             4@\       _       	          @33�?�S����?
             3@]       ^                    @I@      �?             (@������������������������       �                     "@������������������������       �                     @������������������������       �                     @������������������������       �                     �?b       c                    �?և���X�?             @������������������������       �                     @d       e                   �i@      �?             @������������������������       �                     �?������������������������       �                     @g       n                   �l@������?|            `i@h       m                    c@�����?>            @Y@i       j                    �?�����H�?             "@������������������������       �                     @k       l                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        :             W@o       x                    �?l��\��?>            �Y@p       q                    �?�z�G��?             4@������������������������       �                     @r       s                    @I@և���X�?	             ,@������������������������       �                     @t       w                     @؇���X�?             @u       v                   0c@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?y       �                   �t@Ћ����?0            �T@z       {                    �F@ ���J��?-            �S@������������������������       �                     D@|       }                    �?�}�+r��?             C@������������������������       �                     0@~       �                   @[@�C��2(�?             6@       �                   @q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �^@P���Q�?             4@������������������������       �                     $@�       �                     L@ףp=
�?             $@������������������������       �                     @�       �                   p`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   u@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   pb@�&!��?            �E@�       �       	          833�?      �?             A@�       �                    V@z�G�z�?             4@������������������������       �                     @�       �                    �L@�IєX�?             1@������������������������       �        	             (@�       �                   @r@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?@4և���?
             ,@�       �                   pc@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                     "@�       �                    �?@?�8��?�            �w@�       �       
             �?��t����?�            Ps@�       �                   �U@���7�?�            �p@������������������������       �                     �?�       �                    �R@�w�>τ�?�            pp@�       �       
             �?�`�L[,�?�            0p@������������������������       �                     D@�       �                   Pe@���(-�?�            `k@������������������������       �        "             K@�       �                   �Z@�1�`jg�?h            �d@�       �                   a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �D@�@�?f            `d@�       �                   �f@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@�       �                   @a@p�|�i�?_             c@�       �                    �?�T�~~4�?J            @]@�       �                   hu@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�       �                    �?@��!�Q�?B            @Z@������������������������       �        2            �T@�       �                   �_@�nkK�?             7@�       �                   �]@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@�       �                    �?(N:!���?            �A@�       �                    @G@؇���X�?             <@������������������������       �                     �?�       �                    �?�����H�?             ;@�       �                   �a@r�q��?
             2@�       �                    ^@      �?             (@������������������������       �                     @�       �                   `b@      �?              @�       �                    i@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     "@������������������������       �                     @�       �                   �p@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �a@��Hg���?            �F@�       �                   `_@b�h�d.�?            �A@�       �                    �?������?             .@������������������������       �                     @�       �                     N@�8��8��?             (@������������������������       �                      @�       �       	          ����?      �?             @������������������������       �                     �?������������������������       �                     @�       �       	             �?ףp=
�?             4@�       �                   �`@�<ݚ�?             "@������������������������       �                     @�       �                   `k@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                   �]@      �?             $@�       �                    Z@����X�?             @������������������������       �                     �?�       �       	             �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    V@���A��?3            �R@�       �                    �L@      �?             0@������������������������       �                     "@�       �       	          ����?؇���X�?             @������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?П[;U��?%             M@�       �                    �?�I� �?             G@�       �                   `c@>A�F<�?             C@�       �                     N@l��\��?             A@������������������������       �                     6@�       �                    �?      �?             (@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                     N@�8��8��?	             (@������������������������       �                      @�       �       	          ���@      �?             @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�t�b��     h�h(h+K ��h-��R�(KK�KK��h_�B�       �x@     P�@     @u@     `h@     �K@      c@      (@     �X@      (@      I@      &@      6@      @      @               @      @      �?              �?      @              @      3@              ,@      @      @       @      @              @       @              @              �?      <@      �?      "@      �?                      "@              3@             �H@     �E@     �J@      4@      "@      $@      "@       @      "@      @      "@      �?      @              @      �?              @      @      @                      @      @               @              $@              7@      F@      6@      9@      ,@      @      "@              @      @      @      @       @      @       @                      @      @                      @       @      3@      @       @      �?       @      �?                       @       @              @      1@       @      ,@       @                      ,@      @      @      �?      @      �?                      @       @              �?      3@      �?      @              @      �?                      .@     �q@     �E@     0p@      :@      &@      @      @      �?              �?      @               @      @      @              @      @      @                      @      o@      4@     �K@      $@      J@      @     �A@              1@      @      �?       @              �?      �?      �?      �?                      �?      0@      @      0@      @      "@      @      "@                      @      @                      �?      @      @              @      @      �?              �?      @              h@      $@      Y@      �?       @      �?      @              @      �?              �?      @              W@             @W@      "@      ,@      @      @               @      @      @              �?      @      �?      @      �?                      @              �?     �S@      @      S@       @      D@              B@       @      0@              4@       @      �?      �?              �?      �?              3@      �?      $@              "@      �?      @               @      �?              �?       @              @      �?              �?      @              :@      1@      1@      1@      0@      @              @      0@      �?      (@              @      �?      @                      �?      �?      *@      �?       @               @      �?                      &@      "@              L@     pt@      7@     �q@      (@     �o@      �?              &@     �o@      "@     @o@              D@      "@     @j@              K@      "@     �c@      �?      �?              �?      �?               @     `c@       @      "@       @                      "@      @     @b@       @     �\@      �?      &@              &@      �?              �?      Z@             �T@      �?      6@      �?      @              @      �?                      3@      @      ?@      @      8@      �?              @      8@      @      .@      @      "@              @      @      @      �?      @      �?                      @       @                      @              "@              @       @       @               @       @              &@      A@      @      =@      @      &@      @              �?      &@               @      �?      @      �?                      @       @      2@       @      @              @       @      �?              �?       @                      &@      @      @      @       @              �?      @      �?      @                      �?              @     �@@     �D@      �?      .@              "@      �?      @              @      �?      �?      �?                      �?      @@      :@      ?@      .@      ?@      @      ?@      @      6@              "@      @      @      @      @                      @      @                      @               @      �?      &@               @      �?      @      �?       @               @      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJͷ�/hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B88         |       	          ����?n[��L��?C           ��@       ]                    �?`�-��j�?+           �}@       P                    �?H��=6�?�            �x@                          `Q@��`���?�            �t@       
                    �?�eP*L��?            �@@                           �?      �?              @������������������������       �                      @       	                   `_@r�q��?             @������������������������       �                     �?������������������������       �                     @                          �Z@���Q��?             9@������������������������       �                     "@              	             п      �?             0@������������������������       �                     @              	          ����?�eP*L��?	             &@              
             �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     @       +       
             �?(71����?�            �r@       *                   �x@�"U����?!            �I@                           �?(���@��?            �G@                          pe@�X�<ݺ?             2@������������������������       �        	             ,@                          `m@      �?             @������������������������       �                     @������������������������       �                     �?       %                    �?l��[B��?             =@                            �?     ��?	             0@                           �N@���Q��?             @������������������������       �                      @������������������������       �                     @!       $                   �b@�C��2(�?             &@"       #                   pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@&       )                    �O@8�Z$���?
             *@'       (       
             �?�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?������������������������       �                     @,       I       	            �?0��P�?�            �n@-       @                    �?���>4ֵ?�             l@.       ?                   �b@ZՏ�m|�?            �H@/       >                   �_@��E�B��?            �G@0       7                    �?����X�?             5@1       6                   �[@      �?             $@2       3                    �?r�q��?             @������������������������       �                     @4       5                    �H@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @8       9                   �b@�C��2(�?	             &@������������������������       �                     @:       ;                    @I@r�q��?             @������������������������       �                     @<       =                     N@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     :@������������������������       �                      @A       B                    @L@���ib#�?j            �e@������������������������       �        ]             c@C       H                   �m@�C��2(�?             6@D       G                    �?z�G�z�?             $@E       F                   @l@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     (@J       K                   �a@�GN�z�?
             6@������������������������       �                     "@L       M                    �?�n_Y�K�?             *@������������������������       �                     @N       O                   xp@����X�?             @������������������������       �                     @������������������������       �                      @Q       R       
             �?�y(dD�?/            @P@������������������������       �                     B@S       X                   `]@V�a�� �?             =@T       W       	          833�?      �?              @U       V                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @Y       \                   ``@���N8�?             5@Z       [                    V@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �        
             *@^       q                   �b@����[��?8            �S@_       f                   @[@��f/w�?,            �N@`       a                    �D@�8��8��?             8@������������������������       �                     �?b       c       	          ����?�nkK�?             7@������������������������       �                     4@d       e                   p`@�q�q�?             @������������������������       �                      @������������������������       �                     �?g       l       
             �?V������?            �B@h       i                    l@ ��WV�?             :@������������������������       �        
             ,@j       k                   @\@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@m       n                     P@�C��2(�?             &@������������������������       �                     "@o       p       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?r       {                     R@�t����?             1@s       z                    �?z�G�z�?             .@t       u                   @j@      �?             @������������������������       �                      @v       y       	          @33�?      �?             @w       x                    @D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                      @}       �                   �b@4��6_��?           �{@~       �                    �?@�r-��?�             v@       �                    �?H�z�G�?             D@�       �                   �p@�q�q�?             8@�       �                   @l@և���X�?	             ,@�       �                   �`@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@�       �       	          ����?      �?             0@�       �                   �t@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                   �Q@<�jX��?�            �s@�       �                   Pa@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   p`@�-���?�            `s@�       �                    �?p�eU}�?�            �i@�       �                    �R@��w#'�?m            `d@�       �       	          033@p/k%��?l            @d@�       �                     E@p�[&�?_            �a@�       �                   �_@؇���X�?             @������������������������       �                     @�       �                    �?      �?             @�       �                    �C@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �       	          ����? ��ʻ��?Y             a@�       �                   P`@�(\����?7             T@�       �                   Ph@P���Q�?             D@������������������������       �                     8@�       �                     M@      �?             0@�       �                    �?      �?              @�       �                   �^@�q�q�?             @�       �                   l@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     D@������������������������       �        "             L@�       �                    �?�KM�]�?             3@������������������������       �        	             (@�       �                   @X@����X�?             @������������������������       �                     @�       �                   0p@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    �Q@(L���?            �E@�       �                   P`@�#-���?            �A@�       �                   �f@      �?              @�       �                    `@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     ;@�       �       	          033�?      �?              @������������������������       �                     @������������������������       �                     @�       �                   �a@8�Z$���?:             Z@�       �                   @Z@&�a2o��?'            @Q@������������������������       �                     @�       �                   pv@�����D�?%            @P@�       �                    �?     8�?$             P@�       �       
             �?�t����?            �I@�       �       	          ����?�ʈD��?            �E@�       �                   @a@���Q��?             $@�       �                   `^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                    �@@�       �       	          033�?      �?              @������������������������       �                     @�       �                   �\@�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �d@�n_Y�K�?             *@�       �       	             �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                    �A@�       �       	          `ff@��+�ޯ�?:            �V@�       �                    @F@�r*e���?/            �R@������������������������       �        	             (@�       �                    �?V{q֛w�?&             O@�       �       	          ����?      �?             8@�       �                    �J@      �?             $@������������������������       �                     @�       �                   `]@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   0g@@4և���?             ,@�       �                    �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                    �H@�I�w�"�?             C@�       �                    �?�eP*L��?             &@�       �       	          033�?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?�����H�?             ;@�       �                   �p@"pc�
�?	             &@������������������������       �                     @�       �                   `a@����X�?             @������������������������       �                      @������������������������       �                     @�       �                   0d@      �?             0@������������������������       �                     @�       �                    @�����H�?             "@������������������������       �                     @�       �       	          033�?      �?             @������������������������       �                     �?������������������������       �                     @�                           @O@@�0�!��?             1@�       �                    `@��S�ۿ?
             .@������������������������       �                     "@�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KMKK��h_�B       �z@     �~@     `t@     `b@     �r@     �W@     `q@      J@      .@      2@      @      @               @      @      �?              �?      @              $@      .@              "@      $@      @      @              @      @       @      @              @       @              @             pp@      A@      @@      3@      @@      .@      1@      �?      ,@              @      �?      @                      �?      .@      ,@      *@      @      @       @               @      @              $@      �?      �?      �?              �?      �?              "@               @      &@      �?      &@      �?                      &@      �?                      @     �l@      .@     �j@      $@     �D@       @     �D@      @      .@      @      @      @      @      �?      @               @      �?              �?       @                      @      $@      �?      @              @      �?      @               @      �?              �?       @              :@                       @     �e@       @      c@              4@       @       @       @      �?       @      �?                       @      @              (@              1@      @      "@               @      @      @               @      @              @       @              7@      E@              B@      7@      @      @      @      @       @      @                       @              @      4@      �?      @      �?              �?      @              *@              9@     �J@      *@      H@       @      6@      �?              �?      6@              4@      �?       @               @      �?              &@      :@      �?      9@              ,@      �?      &@      �?                      &@      $@      �?      "@              �?      �?              �?      �?              (@      @      (@      @      @      @               @      @      �?       @      �?              �?       @              �?              "@                       @      Z@     Pu@      K@     �r@      7@      1@       @      0@       @      @       @      @       @                      @      @                      $@      .@      �?      @      �?      @                      �?      $@              ?@     �q@      @      �?      @                      �?      <@     �q@      (@     @h@      @     �c@      @     �c@      @     �a@      �?      @              @      �?      @      �?       @               @      �?                      �?       @     �`@       @     �S@       @      C@              8@       @      ,@       @      @       @      @      �?      @      �?                      @      �?                       @               @              D@              L@       @      1@              (@       @      @              @       @       @               @       @              �?              @     �B@      @      @@      @      @      �?      @              @      �?               @                      ;@      @      @      @                      @      0@      V@      0@     �J@      @              (@     �J@      &@     �J@      @     �F@      @     �C@      @      @      @      �?              �?      @                      @             �@@       @      @              @       @      �?      �?      �?      �?                      �?      �?              @       @       @       @       @                       @      @              �?                     �A@      I@     �D@     �G@      ;@      (@             �A@      ;@      @      2@      @      @              @      @      �?              �?      @              �?      *@      �?      �?      �?                      �?              (@      =@      "@      @      @      @      @              @      @                      @      8@      @      "@       @      @              @       @               @      @              .@      �?      @               @      �?      @              @      �?              �?      @              @      ,@      �?      ,@              "@      �?      @              @      �?               @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ%�}+hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKh~�BH4         z                    �?���3L�?:           ��@       G       
             �?��b��?<           H�@       
                    b@�8��8��?�            �x@              	          ����?�Ń��̧?D            �_@������������������������       �        7             Y@       	       
             �?ȵHPS!�?             :@                           �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �        
             4@                          �Q@�����H�?�            �p@������������������������       �                     �?       2       	          pff�? �ߙ���?�            �p@                           �?|��+�?^            �b@                          �f@�q�q�?             ;@������������������������       �                     @                          �^@      �?             8@������������������������       �                      @                          hu@"pc�
�?             6@                           �G@ףp=
�?             4@������������������������       �                      @������������������������       �        	             2@������������������������       �                      @                          �e@�R����?N            @^@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                           �?U���y�?L            �]@������������������������       �                     4@              	          ����?�����H�?>            �X@������������������������       �                     @@        %                    @L@� y���?,            �P@!       $       	          ����?P���Q�?             D@"       #                    �?�����H�?             2@������������������������       �                      @������������������������       �                     0@������������������������       �                     6@&       )                    �L@�q�q�?             ;@'       (                   n@����X�?             @������������������������       �                     @������������������������       �                      @*       /                   �b@z�G�z�?             4@+       ,                   �o@�t����?             1@������������������������       �        	             (@-       .                   p`@���Q��?             @������������������������       �                      @������������������������       �                     @0       1                    �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?3       F                    �R@0 �����?I            @^@4       5                   �Z@Xc!J�ƴ?H            �]@������������������������       �                     �?6       =       	          033@ȑ����?G            @]@7       8                    c@ ��PUp�?.            �Q@������������������������       �        +            �P@9       :                    _@      �?             @������������������������       �                      @;       <                    q@      �?              @������������������������       �                     �?������������������������       �                     �?>       ?                   8p@���.�6�?             G@������������������������       �                     ;@@       E                    `@�S����?             3@A       B       
             �?      �?              @������������������������       �                     @C       D                   �^@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     &@������������������������       �                     @H       [                    P@l��TO��?P            @_@I       V                   �`@tk~X��?             B@J       Q                    �?����X�?             5@K       P       	          `ff�?�r����?	             .@L       O       	          ����?@4և���?             ,@M       N                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?R       U                   �a@�q�q�?             @S       T                   `[@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @W       Z                    �?��S�ۿ?             .@X       Y                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@\       s                    �?:��?:            @V@]       b                   �a@��d��?*            �O@^       _                   p@      �?             @@������������������������       �                     :@`       a       	             �?r�q��?             @������������������������       �                     @������������������������       �                     �?c       l                     N@¦	^_�?             ?@d       k                    @J@�<ݚ�?             ;@e       h                   �e@�z�G��?             4@f       g                   @_@d}h���?	             ,@������������������������       �                     @������������������������       �                     &@i       j                   l@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @m       r       	          @33�?      �?             @n       o                   �i@�q�q�?             @������������������������       �                     �?p       q                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?t       u                   �a@�θ�?             :@������������������������       �                     0@v       w                   @b@���Q��?             $@������������������������       �                     @x       y                   �_@�q�q�?             @������������������������       �                     @������������������������       �                      @{       �                    �K@Z��m��?�            �x@|       �       	          033�? ���$�?�            �o@}       �                   �c@�����?�            �l@~       �       	             �?���Q��?             .@       �                    @C@      �?	             (@������������������������       �                     @�       �                    �?�q�q�?             "@�       �                    �?r�q��?             @�       �                   �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   @`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?p)�����?�             k@������������������������       �        N            �_@�       �                    @K@ ��~���?<            �V@�       �                   �n@�t����?8            @U@�       �                   �c@�g�y��?'             O@�       �                   �l@0�)AU��?#            �L@������������������������       �                     C@�       �                   @m@�}�+r��?             3@�       �                   `e@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             ,@�       �       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?�LQ�1	�?             7@�       �                    �?�q�q�?             (@������������������������       �                      @�       �                    �I@z�G�z�?             $@������������������������       �                     @�       �                   �r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             &@�       �       
             �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    �?�û��|�?             7@�       �       
             �?����X�?             @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    m@      �?
             0@�       �                    �J@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�       �                   (p@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   �b@l���?\            �a@�       �       
             �?�q�Q�??             X@�       �       
             �?��X���?-            @Q@�       �                   a@�q�q�?             @�       �                   @]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   b@؇���X�?(            �O@�       �                    �O@�3Ea�$�?              G@�       �                   �^@��� ��?             ?@�       �                   �^@ �q�q�?             8@�       �                    @M@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@�       �       	          ����?և���X�?             @������������������������       �                      @�       �                    �?���Q��?             @������������������������       �                     �?�       �                   �`@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?�q�q�?	             .@�       �                     Q@����X�?             @�       �                   �_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     1@�       �                   �a@�����H�?             ;@������������������������       �                     5@�       �                    �?      �?             @������������������������       �                     �?�       �                   �b@���Q��?             @������������������������       �                      @�       �                   �Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   0d@��[�p�?            �G@�       �                    @HP�s��?             9@������������������������       �                     5@�       �                   `c@      �?             @������������������������       �                      @������������������������       �                      @�       �                    @L@���|���?             6@������������������������       �                     @�       �                    b@��.k���?             1@�       �                   @_@      �?              @�       �                    ]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�<ݚ�?             "@�       �                    c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       px@     x�@     �X@     `z@     �@@     �v@      @     �^@              Y@      @      7@      @      @      @                      @              4@      >@      n@      �?              =@      n@      5@     �_@      "@      2@      @              @      2@       @              @      2@       @      2@       @                      2@       @              (@     @[@      �?      �?      �?                      �?      &@      [@              4@      &@      V@              @@      &@      L@       @      C@       @      0@       @                      0@              6@      "@      2@      @       @      @                       @      @      0@       @      .@              (@       @      @       @                      @       @      �?       @                      �?       @     @\@      @     @\@      �?              @     @\@      �?     �Q@             �P@      �?      @               @      �?      �?              �?      �?              @     �E@              ;@      @      0@      @      @              @      @       @               @      @                      &@      @             �P@     �M@      @      =@      @      .@       @      *@      �?      *@      �?      �?      �?                      �?              (@      �?              @       @      �?       @      �?                       @      @              �?      ,@      �?      �?      �?                      �?              *@     �M@      >@     �J@      $@      ?@      �?      :@              @      �?      @                      �?      6@      "@      5@      @      ,@      @      &@      @              @      &@              @      @              @      @              @              �?      @      �?       @              �?      �?      �?      �?                      �?              �?      @      4@              0@      @      @      @               @      @              @       @             @r@     @Z@     @k@      B@      j@      6@      @      "@      @      @              @      @      @      @      �?      �?      �?              �?      �?              @              �?       @               @      �?                      @     `i@      *@     �_@             @S@      *@     �R@      $@      N@       @      L@      �?      C@              2@      �?      @      �?              �?      @              ,@              @      �?      @                      �?      .@       @      @       @       @               @       @              @       @      �?              �?       @              &@               @      @              @       @              "@      ,@      @       @       @       @       @                       @      @              @      (@      �?      &@              &@      �?              @      �?      @                      �?     �R@     @Q@     �B@     �M@      *@      L@      @       @      �?       @      �?                       @      @              "@      K@      "@     �B@      @      ;@      �?      7@      �?      @      �?                      @              2@      @      @               @      @       @              �?      @      �?      �?      �?      �?                      �?       @              @      $@      @       @       @       @       @                       @      @                       @              1@      8@      @      5@              @      @      �?               @      @               @       @      �?              �?       @             �B@      $@      7@       @      5@               @       @       @                       @      ,@       @      @              "@       @       @      @       @      �?              �?       @                      @      @       @      �?       @      �?                       @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�BH;         �                    �?n[��L��?E           ��@       [       
             �?�)�0z�?:           @                          `_@��u}���?�            Pv@                           �Q@��4+̰�?z            @h@              	          `ff@`Ql�R�?t            �g@                          ``@`��>�ϗ?g            @e@                           @L@�g<a�?1            @S@������������������������       �                     E@	       
                    �? >�֕�?            �A@������������������������       �                     0@                           �L@�KM�]�?             3@������������������������       �                     �?                          �_@�X�<ݺ?             2@������������������������       �        	             ,@                          p`@      �?             @������������������������       �                      @              	          433�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        6            @W@                          �_@�����H�?             2@                          �\@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        
             ,@                           �?�q�q�?             @������������������������       �                     �?                          �p@z�G�z�?             @������������������������       �                     @������������������������       �                     �?       8                    �?X�Բ���?j            `d@        !                    `@���!pc�?            �@@������������������������       �                     �?"       )       	          hff�?      �?             @@#       (                    �?�q�q�?             @$       '                    �?z�G�z�?             @%       &       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?*       7                    �?8�Z$���?             :@+       2                   pl@�㙢�c�?             7@,       -                   �`@      �?             @������������������������       �                     �?.       1                   �a@���Q��?             @/       0       	             �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?3       6       	          ����?�IєX�?             1@4       5                   �u@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     @9       :       	          833�?���Ls�?R            @`@������������������������       �                     ?@;       D                   `@<���D�??            �X@<       C                   l@�����?
             3@=       B                    �?      �?             (@>       ?                    �F@�q�q�?             "@������������������������       �                      @@       A                    @K@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @E       J                   pb@��(\���?5             T@F       I                    �?���J��?"            �I@G       H                    �J@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     F@K       N                   �b@д>��C�?             =@L       M                   l@      �?             @������������������������       �                     @������������������������       �                     @O       P       
             �?���}<S�?             7@������������������������       �                     @Q       Z                   `c@�����H�?             2@R       Y                   0c@"pc�
�?             &@S       T                   �q@ףp=
�?             $@������������������������       �                     @U       X                   �b@      �?             @V       W                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @\       �                    �?N� ˔x�?V            �a@]       z                    �?���vq�?B            �Z@^       o                    @N@�P�����?0            �S@_       n       	          ����?pH����?)            �P@`       i                    @F@X��Oԣ�?'             O@a       b                   �b@�θ�?             :@������������������������       �                     "@c       d                    �?ҳ�wY;�?	             1@������������������������       �                     @e       f                   pf@8�Z$���?             *@������������������������       �                     $@g       h                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?j       k                    �?������?             B@������������������������       �                      @l       m                   @E@h�����?             <@������������������������       �                     �?������������������������       �                     ;@������������������������       �                     @p       w       	          ����?      �?             (@q       r                   �i@����X�?             @������������������������       �                     @s       v                    �?�q�q�?             @t       u                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?x       y                    ]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @{       �       	             �?������?             ;@|       �                   �a@��
ц��?	             *@}       ~                    h@�<ݚ�?             "@������������������������       �                     @       �                   �r@���Q��?             @�       �                   �`@�q�q�?             @������������������������       �                     �?�       �                     G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?@4և���?	             ,@������������������������       �                      @�       �                    c@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �`@@�0�!��?             A@�       �                   �Y@�8��8��?             8@������������������������       �                     �?�       �                    ]@�nkK�?             7@������������������������       �                     4@�       �                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    b@���Q��?             $@�       �                   �a@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �K@���CZ��?           Pz@�       �                    �?4hy���?�            �q@�       �       
             �?�*0��
�?�            `o@�       �                   �f@#z�i��?            �D@�       �                    �G@�<ݚ�?             "@�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �a@     ��?             @@�       �                    �?      �?             @�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �       	          ���@؇���X�?             <@�       �                    �?�����H�?             ;@�       �                    �?$�q-�?             :@������������������������       �                     5@�       �                    �H@���Q��?             @�       �                   �_@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �?P�c0"�?�            @j@�       �                    �?ܷ��?��?             =@������������������������       �                     ,@�       �                   �b@z�G�z�?	             .@������������������������       �                      @�       �                   xp@$�q-�?             *@������������������������       �                     &@�       �                   xr@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?@�:;��?q            �f@�       �                   @n@@=��?`            �c@������������������������       �        7            �W@�       �                   �n@     ��?)             P@������������������������       �                     �?������������������������       �        (            �O@������������������������       �                     7@�       �                    I@)O���?             B@������������������������       �                     @�       �       
             �?`՟�G��?             ?@�       �                     J@��S�ۿ?             .@������������������������       �                     &@�       �                   �`@      �?             @������������������������       �                      @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@�       �                    �?��:c���?W            �`@�       �                    �?�n_Y�K�?=            �V@�       �                    �?��f/w�?*            �N@�       �                    ]@��>4և�?             <@������������������������       �                     �?�       �                    �?��}*_��?             ;@�       �                   �l@�q�q�?             @������������������������       �                     �?�       �                    @L@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �       	          033�?����X�?             5@�       �                    q@@�0�!��?             1@������������������������       �                     (@�       �                    c@���Q��?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   m@�FVQ&�?            �@@������������������������       �        
             *@�       �       
             �?ףp=
�?             4@�       �                   �_@      �?             @�       �                   8p@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@�       �       	          @33�?������?             >@������������������������       �                     &@�       �       	          ����?D�n�3�?             3@������������������������       �                     @�       �                    �N@     ��?             0@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    �?z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �[@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�                          �?�K��&�?            �E@�       �                   a@      �?             (@������������������������       �                     @                         Pc@      �?             @������������������������       �                     @������������������������       �                     @                        �`@¦	^_�?             ?@������������������������       �        
             1@            	             �?X�Cc�?	             ,@������������������������       �                     @            	             �?X�<ݚ�?             "@������������������������       �                      @	                          P@և���X�?             @
                        `^@z�G�z�?             @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KMKK��h_�B�       �z@     �~@     �Z@     px@      ;@     �t@      @     �g@      @      g@       @      e@       @     �R@              E@       @     �@@              0@       @      1@      �?              �?      1@              ,@      �?      @               @      �?      �?      �?                      �?             @W@       @      0@       @       @       @                       @              ,@       @      @      �?              �?      @              @      �?              5@     �a@      "@      8@      �?               @      8@      @       @      @      �?      �?      �?              �?      �?              @                      �?      @      6@      @      3@      @      @      �?               @      @       @       @               @       @                      �?      �?      0@      �?      @              @      �?                      "@              @      (@     �]@              ?@      (@     �U@      @      *@      @      @      @      @       @              �?      @              @      �?              @                      @      @     �R@      �?      I@      �?      @      �?                      @              F@      @      8@      @      @      @                      @       @      5@              @       @      0@       @      "@      �?      "@              @      �?      @      �?      �?              �?      �?                       @      �?                      @     �S@     �N@     @R@     �@@     �P@      *@      N@      @     �K@      @      4@      @      "@              &@      @              @      &@       @      $@              �?       @               @      �?             �A@      �?       @              ;@      �?              �?      ;@              @              @      @       @      @              @       @      �?      �?      �?              �?      �?              �?              @      �?              �?      @              @      4@      @      @       @      @              @       @      @       @      �?      �?              �?      �?              �?      �?                       @      @              �?      *@               @      �?      @              @      �?              @      <@       @      6@      �?              �?      6@              4@      �?       @      �?                       @      @      @      @      @      @                      @              @     @t@     @X@     @o@     �B@      m@      2@      ;@      ,@       @      @       @      �?       @                      �?              @      9@      @      �?      @      �?      �?      �?                      �?               @      8@      @      8@      @      8@       @      5@              @       @      �?       @      �?                       @       @                      �?              �?     �i@      @      :@      @      ,@              (@      @               @      (@      �?      &@              �?      �?              �?      �?             �f@      �?     �c@      �?     �W@             �O@      �?              �?     �O@              7@              1@      3@              @      1@      ,@      �?      ,@              &@      �?      @               @      �?      �?              �?      �?              0@             �R@      N@      L@     �A@      H@      *@      1@      &@              �?      1@      $@       @      @      �?              �?      @      �?                      @      .@      @      ,@      @      (@               @      @      �?              �?      @      �?                      @      �?      @              @      �?              ?@       @      *@              2@       @       @       @       @      �?       @                      �?              �?      0@               @      6@              &@       @      &@      @              @      &@      @       @              �?      @      �?      @              �?      �?              �?      �?              �?      "@      �?                      "@      2@      9@      "@      @      @              @      @              @      @              "@      6@              1@      "@      @      @              @      @               @      @      @      @      �?      �?      �?              �?      �?              @                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��iXhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK煔h~�B�2         .                    _@�&���?Q           ��@              
             �?zI�^�p�?u             g@                           �?������?S             a@       	                    �Q@`'�J�?@            �Y@                          `X@�q�q�?=             X@                           X@�}�+r��?             3@������������������������       �        
             2@������������������������       �                     �?������������������������       �        2            @S@
                          @L@      �?             @������������������������       �                     @������������������������       �                     @              	             @H�V�e��?             A@                          �]@�r����?             >@������������������������       �        	             0@                           �?����X�?             ,@                            K@և���X�?             @������������������������       �                      @              
             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @                            L@      �?             @������������������������       �                     �?������������������������       �                     @       '                    �?���Q �?"            �H@       &                   @E@      �?             @@                          �]@��a�n`�?             ?@              	          ����?և���X�?             @������������������������       �                     @������������������������       �                     @        !                    �M@      �?             8@������������������������       �                     3@"       #       	             �?���Q��?             @������������������������       �                     �?$       %                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?(       -                    �?��.k���?             1@)       ,       	          ����?�	j*D�?	             *@*       +                   �b@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @������������������������       �                      @������������������������       �                     @/       �       
             �?\Ǒ��?�           �@0       s                   �`@B@!�S3�?�            0x@1       R                    �?�j&|mH�?�            @h@2       ;                    �?�w��d��??            @W@3       :                    �?z�G�z�?             9@4       5                   `X@�LQ�1	�?             7@������������������������       �                     �?6       9                    �?�C��2(�?             6@7       8       	          ����?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     (@������������������������       �                      @<       E       	          ����?��paR�?.             Q@=       B                   �`@؇���X�?             <@>       A                    �? �q�q�?             8@?       @       
             �?�}�+r��?             3@������������������������       �                     �?������������������������       �                     2@������������������������       �                     @C       D                   �u@      �?             @������������������������       �                     @������������������������       �                     �?F       G                    ]@H�z�G�?             D@������������������������       �                      @H       Q                     P@     ��?             @@I       J       	          ����?��>4և�?             <@������������������������       �                     *@K       P                    @������?             .@L       M                    �?d}h���?             ,@������������������������       �        	             $@N       O                    �L@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @S       r                    �?L��/�/�?D            @Y@T       U                   �Y@̘SJl��?7            �S@������������������������       �        	             .@V       [                   `\@     ��?.             P@W       Z                   @q@      �?             $@X       Y                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @\       e                   �\@�+$�jP�?)             K@]       ^                    �?���Q��?	             $@������������������������       �                      @_       `       	          ����?      �?              @������������������������       �                      @a       b                     M@�q�q�?             @������������������������       �                     @c       d                    l@�q�q�?             @������������������������       �                     �?������������������������       �                      @f       m                   �b@�C��2(�?              F@g       l       	          ����?�}�+r��?             C@h       i                   �q@�<ݚ�?             "@������������������������       �                     @j       k                     K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     =@n       o                    �?�q�q�?             @������������������������       �                      @p       q                   `e@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     6@t       �                   �b@�׾���?x             h@u       �                    �?��<�Ұ?]            `b@v       {                    �?�T�~~4�?L            @]@w       z       	             �?�X�<ݺ?             2@x       y                    �J@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@|       �                   �[@`�LVXz�?@            �X@}       �                   �a@�X�<ݺ?             2@~                           g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@������������������������       �        2            @T@�       �                   pb@ףp=
�?             >@������������������������       �                     8@�       �       	             �?      �?             @������������������������       �                      @�       �                   `c@      �?             @������������������������       �                      @�       �                    e@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `a@�I� �?             G@������������������������       �                     @�       �                    �?���?            �D@�       �                    �?�LQ�1	�?             7@�       �                   �b@�eP*L��?             &@������������������������       �                     @������������������������       �                     @�       �       	          pff�?      �?             (@������������������������       �                     �?�       �                    @"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�       �                   hr@�����H�?             2@������������������������       �        	             ,@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?E�Vl��?�            �u@�       �                   �k@`�H{�i�?�            s@�       �                    �?Pa�	�?\            �`@�       �                    f@�����?             5@������������������������       �                     �?�       �                     G@P���Q�?             4@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@�       �                    @N@�Μ�5�?P            �[@�       �                    �?@�n���?I            �Y@�       �                    �I@�a�O�?D            @X@������������������������       �        ,             O@�       �                   �_@��?^�k�?            �A@�       �                    �?�8��8��?             (@�       �                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     7@������������������������       �                     @�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    �?��	= ��?k            �e@�       �                    �M@������?            �F@�       �                    �L@� ��1�?            �D@�       �                    �?��hJ,�?             A@�       �                   �c@�q�q�?             "@�       �                    ^@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    ]@HP�s��?             9@�       �       	          ����?      �?              @�       �                    �H@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     1@�       �                   p`@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �L@     8�?M             `@������������������������       �        ;            �X@�       �                   �s@r�q��?             >@�       �                    �?�����H�?             ;@�       �                    m@���7�?             6@������������������������       �                     �?������������������������       �                     5@�       �                   �_@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �e@#z�i��?            �D@�       �                    �?      �?             B@�       �                    �?��� ��?             ?@�       �       	          ����?��2(&�?             6@�       �                   @`@�z�G��?             $@������������������������       �                     @�       �                    a@      �?             @������������������������       �                      @�       �                    d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                    �G@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�t�b��     h�h(h+K ��h-��R�(KK�KK��h_�Bp        y@      �@      <@     �c@      &@     @_@      @     �X@      �?     �W@      �?      2@              2@      �?                     @S@      @      @      @                      @      @      ;@      @      :@              0@      @      $@      @      @       @               @      @       @                      @              @      @      �?              �?      @              1@      @@       @      8@      @      8@      @      @      @                      @      @      5@              3@      @       @              �?      @      �?      @                      �?      �?              "@       @      "@      @      "@       @      "@                       @               @              @     `w@     pv@      S@     ps@      L@     @a@     �D@      J@      4@      @      4@      @              �?      4@       @       @       @               @       @              (@                       @      5@     �G@      @      8@      �?      7@      �?      2@      �?                      2@              @      @      �?      @                      �?      1@      7@               @      1@      .@      1@      &@      *@              @      &@      @      &@              $@      @      �?      @                      �?      �?                      @      .@     �U@      .@      P@              .@      .@     �H@      @      @      @      �?              �?      @                      @      $@      F@      @      @               @      @       @       @              @       @      @              �?       @      �?                       @      @      D@       @      B@       @      @              @       @      �?              �?       @                      =@       @      @               @       @       @       @                       @              6@      4@     �e@      @     �a@       @     �\@      �?      1@      �?      @      �?                      @              &@      �?     �X@      �?      1@      �?      �?              �?      �?                      0@             @T@      @      ;@              8@      @      @               @      @      �?       @              �?      �?              �?      �?              .@      ?@      @              $@      ?@       @      .@      @      @      @                      @      @      "@      �?               @      "@              "@       @               @      0@              ,@       @       @       @                       @     �r@      H@     �q@      5@      `@      @      3@       @              �?      3@      �?      @      �?              �?      @              .@             @[@       @     �Y@      �?      X@      �?      O@              A@      �?      &@      �?      �?      �?              �?      �?              $@              7@              @              @      �?              �?      @             �c@      1@     �@@      (@     �@@       @      =@      @      @      @       @      @       @                      @      @              7@       @      @       @      @       @      @                       @       @              1@              @      @              @      @                      @     �^@      @     �X@              9@      @      8@      @      5@      �?              �?      5@              @       @               @      @              �?       @               @      �?              ,@      ;@      "@      ;@      @      ;@      @      3@      @      @              @      @      �?       @              �?      �?              �?      �?                      (@      �?       @      �?                       @      @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�1\ hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �                    �?\r��ۖ�?[           ��@       K       
             �?��#>֍�?X           �@       "                    �?@��C�?z            `f@                          �n@HP�s��?F             Y@                          P`@������?/             R@������������������������       �                     H@              	          ����?�8��8��?             8@              	            �?8�Z$���?             *@	                          �b@�8��8��?
             (@
                          �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?������������������������       �                     &@                          �Q@d}h���?             <@������������������������       �                     �?       !                   �e@�+$�jP�?             ;@                           �?8�Z$���?             :@              	          ����?և���X�?             @                           �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                          Pr@�}�+r��?             3@������������������������       �                     $@                           �?�����H�?             "@������������������������       �                     �?              	             �?      �?              @������������������������       �                     @                            �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?#       0                    �?bf@����?4            �S@$       /                    �?�C��2(�?             6@%       *                    @L@ףp=
�?             4@&       )                     H@��S�ۿ?             .@'       (                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @+       .                    �?z�G�z�?             @,       -                   �j@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @1       >                   0a@���b���?%            �L@2       =                    @L@�eP*L��?            �@@3       <                   hp@ �o_��?             9@4       ;                   @W@"pc�
�?             6@5       :                    @�q�q�?             @6       9                    �?      �?             @7       8                    @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     0@������������������������       �                     @������������������������       �                      @?       B                    �J@�q�q�?             8@@       A                    �?      �?             @������������������������       �                      @������������������������       �                      @C       J       	          ���@R���Q�?             4@D       I                    W@�X�<ݺ?             2@E       H                    �?r�q��?             @F       G                     P@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             (@������������������������       �                      @L       U                    �?������?�             u@M       N                   s@г�wY;�?B            �Y@������������������������       �        5            @U@O       T                    �?@�0�!��?             1@P       S                   �b@���Q��?             @Q       R                    @L@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     (@V       �                    �?:�&���?�            @m@W       p                    �?pLBQh��?�             i@X       ]                    �?x��}�?$            �K@Y       Z                   �a@      �?             $@������������������������       �                     @[       \                   @^@����X�?             @������������������������       �                     @������������������������       �                      @^       c                   @E@:	��ʵ�?            �F@_       `       	          @33�?      �?             @������������������������       �                     �?a       b                    a@�q�q�?             @������������������������       �                      @������������������������       �                     �?d       o                    �?�p ��?            �D@e       n                    b@V�a�� �?             =@f       m                    �N@ȵHPS!�?             :@g       h                    @I@ �q�q�?             8@������������������������       �                     0@i       l       	          @33�?      �?              @j       k                    @J@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     (@q       �                    �?�F��O�?^            @b@r       �                   �c@����X�?             5@s       |       	          ����?���y4F�?             3@t       {                   �d@��S�ۿ?	             .@u       z       	          @33�?؇���X�?             @v       w                   Pl@r�q��?             @������������������������       �                     @x       y                    �O@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @}       ~                   0b@      �?             @������������������������       �                      @       �                    e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �O@H�Swe�?P            @_@�       �                   @[@��7�K¨?N            @^@�       �                    �G@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   @p@�T�~~4�?J            @]@������������������������       �        6             U@�       �                   Xp@�FVQ&�?            �@@������������������������       �                      @������������������������       �                     ?@�       �                   Pc@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�'�=z��?            �@@�       �                   @[@�E��ӭ�?             2@������������������������       �        	             *@������������������������       �                     @�       �       	          ����?������?             .@������������������������       �        	             $@�       �                   �Z@z�G�z�?             @������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �J@�חF�P�?           0y@�       �                   Hq@� Mv:�?\            �`@�       �                   �b@�{���2�?I            �[@�       �                   �a@��wy���?;             W@�       �       
             �?      �?0             R@�       �                   �U@�U�=���?+            �P@������������������������       �                      @�       �                    �?     �?*             P@�       �       	          pff�?@3����?$             K@������������������������       �                     =@�       �       	          ����?`2U0*��?             9@������������������������       �                     �?������������������������       �                     8@�       �                    �I@z�G�z�?             $@�       �       
             �?�����H�?             "@������������������������       �                     @�       �                     H@r�q��?             @�       �                    �F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    I@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   `c@      �?             4@�       �                    �?����X�?             ,@�       �                   @Z@r�q��?             (@������������������������       �                      @������������������������       �                     $@������������������������       �                      @������������������������       �                     @�       �                    �I@���y4F�?             3@�       �                    V@�t����?             1@������������������������       �                     �?�       �       
             �?      �?             0@�       �                    @C@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     8@�       �       	          ����?T�P*�/�?�            �p@�       �       
             �?$gv&��?G            �]@�       �                   �_@������?8            @X@�       �                   �Z@���N8�?             5@�       �                   �p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     2@�       �                   Pn@$�Z����?+             S@�       �                    �K@�&=�w��?            �J@�       �                    Y@�q�q�?             @������������������������       �                     @�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �G@�       �                     N@�û��|�?             7@�       �                    �?�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �       	          ����?և���X�?             ,@������������������������       �                     @�       �                   �p@z�G�z�?             $@������������������������       �                     @�       �                   `]@      �?             @������������������������       �                     �?�       �                    @O@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    h@և���X�?             5@������������������������       �                     @�       �                    �?�t����?             1@�       �                   �d@X�<ݚ�?             "@�       �       	          ����?r�q��?             @�       �                   Pa@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�                          @�U�e?Ƕ?`            �b@�                          @N@xL��N�?^            �b@�       �                   �b@�>����?2            @T@�       �                   0i@�kb97�?0            @S@�       �       	             �?�㙢�c�?             7@�       �                    �?      �?              @�       �                    �K@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?��S�ۿ?
             .@�       �                    @M@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        "             K@�                          �c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        ,            �P@                         �?      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KMKK��h_�BP       py@     �@     `u@     �e@     �I@      `@       @      W@       @     �Q@              H@       @      6@       @      &@      �?      &@      �?       @               @      �?                      "@      �?                      &@      @      6@      �?              @      6@      @      6@      @      @      @      �?      @                      �?              @      �?      2@              $@      �?       @              �?      �?      @              @      �?      �?      �?                      �?      �?             �E@      B@      4@       @      2@       @      ,@      �?      @      �?      @                      �?       @              @      �?       @      �?       @                      �?       @               @              7@      A@      2@      .@      2@      @      2@      @       @      @       @       @      �?       @               @      �?              �?                       @      0@                      @               @      @      3@       @       @               @       @              @      1@      �?      1@      �?      @      �?      @              @      �?                      �?              (@       @             0r@     �F@     �X@      @     @U@              ,@      @       @      @       @       @       @                       @              �?      (@              h@      E@      f@      9@      E@      *@      @      @      @               @      @              @       @             �B@       @       @       @      �?              �?       @               @      �?             �A@      @      7@      @      7@      @      7@      �?      0@              @      �?      @      �?              �?      @               @                       @              @      (@             �`@      (@      .@      @      .@      @      ,@      �?      @      �?      @      �?      @               @      �?              �?       @              �?               @              �?      @               @      �?      �?      �?                      �?               @     �]@      @     �]@      @      @      �?      �?      �?      �?                      �?       @             �\@       @      U@              ?@       @               @      ?@              �?      @      �?                      @      0@      1@      @      *@              *@      @              &@      @      $@              �?      @              @      �?      �?              �?      �?             @P@      u@      A@     @Y@      A@     @S@      3@     @R@      "@     �O@      @     �N@       @              @     �N@      �?     �J@              =@      �?      8@      �?                      8@       @       @      �?       @              @      �?      @      �?       @               @      �?                      @      �?              @       @               @      @              $@      $@      $@      @      $@       @               @      $@                       @              @      .@      @      .@       @              �?      .@      �?      @      �?              �?      @               @                       @              8@      ?@     �m@      8@     �W@      (@     @U@      �?      4@      �?       @      �?                       @              2@      &@     @P@       @     �I@       @      @              @       @      �?              �?       @                     �G@      "@      ,@      �?       @               @      �?               @      @              @       @       @      @               @       @              �?       @      �?       @                      �?      (@      "@              @      (@      @      @      @      �?      @      �?      �?      �?                      �?              @      @               @              @     �a@      @     �a@      @     �R@      @     @R@      @      3@      @      @      @      �?              �?      @                      @      �?      ,@      �?      @              @      �?                      @              K@       @       @       @                       @             �P@      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�5         �       
             �?n�A��?;           ��@       s                   �b@��G���?B           0�@                           �?���AS��?           @{@                           �?JJ����?            �G@              	          ����?�θ�?             :@                          �Z@�q�q�?             @������������������������       �                     �?       	                    �?z�G�z�?             @������������������������       �                     @
                           f@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?ףp=
�?             4@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?                          Po@�X�<ݺ?             2@                          `a@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@                           �?���N8�?
             5@                           @N@�IєX�?             1@������������������������       �                     (@              	          pff�?z�G�z�?             @������������������������       �                     @                          �m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       0                   �[@�̻`mk�?�            Px@        !                   `_@ \� ���?            �H@������������������������       �                     3@"       /                    �?���Q��?             >@#       $                     E@�q�����?             9@������������������������       �                     @%       &                   �Z@p�ݯ��?
             3@������������������������       �                     @'       .                    �?      �?             ,@(       )                   �`@��
ц��?             *@������������������������       �                     @*       -                   �m@؇���X�?             @+       ,       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @1       n                   `f@�q�Y��?�            @u@2       3                   �Q@X(r ԟ�?�            �t@������������������������       �                     �?4       S                    �?���>+T�?�            �t@5       R                   Pp@���2j��?:            �Y@6       G                   �a@,sI�v�?4            �V@7       F                    �?t�e�í�?&            �P@8       E                    `Q@4?,R��?             B@9       >                   �X@(N:!���?            �A@:       =                   �]@�q�q�?             @;       <                   @`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @?       @       
             �? 	��p�?             =@������������������������       �                     �?A       B                   �`@h�����?             <@������������������������       �        	             .@C       D                   �a@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?������������������������       �                     ?@H       Q                    p@��+7��?             7@I       J                   `g@R���Q�?             4@������������������������       �                     $@K       P                    @N@�z�G��?             $@L       O                    �L@���Q��?             @M       N                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     (@T       [       
             �?@�?1X�?�            �l@U       Z                   �\@ףp=
�?             >@V       Y       	             @�θ�?	             *@W       X                    �R@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     1@\       i                    a@�ʱ�O+�?�            �h@]       h       	          ����?�h%�M��?p            `e@^       _       	          ����?      �?,             P@������������������������       �                     >@`       a                    �K@�IєX�?             A@������������������������       �                     ,@b       c       	          hff�?ףp=
�?             4@������������������������       �                     �?d       g                   `X@�}�+r��?             3@e       f                   �W@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             0@������������������������       �        D            �Z@j       k                   pb@@4և���?             <@������������������������       �                     3@l       m                     M@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @o       r                    a@      �?              @p       q                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @t       �                   �b@�p ��?2            �T@u       �       	          ����?� �	��?.            �R@v       {                    �?z�G�z�?             4@w       z                    �?���Q��?             @x       y                   `d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @|       }                   �`@��S�ۿ?	             .@������������������������       �                     *@~                          �d@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�2�o�U�?!            �K@�       �                    �?և���X�?             <@�       �                   �c@���Q��?             4@�       �       	          `ff�?�����H�?             "@������������������������       �                     @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   Po@���|���?             &@�       �                    ^@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �e@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �? 7���B�?             ;@������������������������       �                     6@�       �                    �?z�G�z�?             @������������������������       �                     @�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    @L@ڬ�\mE�?�             y@�       �       	          ����?lI*Lݮ�?�            �q@�       �                    �?Pq�����?�            �o@�       �                   i@�r����?             >@�       �                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @e@ �Cc}�?             <@�       �                    _@�>����?             ;@�       �                    �?�q�q�?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     5@������������������������       �                     �?�       �                    I@���
���?�             l@�       �                    �?և���X�?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	          ����?����q�?�            @k@�       �                   �k@�)ȫ���?}             i@������������������������       �        9            @X@�       �                   �b@ ��WV�?D             Z@������������������������       �                    �I@�       �                    c@�NW���?&            �J@������������������������       �                      @�       �                    l@`'�J�?%            �I@�       �                    b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   0d@��<b�ƥ?"             G@�       �                    �?@4և���?             ,@������������������������       �        
             (@�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @@������������������������       �                     1@�       �                   `U@|��?���?             ;@������������������������       �                     "@�       �       	          ����?�<ݚ�?             2@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             *@�       �       	          pff�?��Q:��?@            �]@�       �                    �M@�G�z.�?+             T@�       �                    �?��
ц��?             :@�       �                   `b@�z�G��?             $@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   `]@     ��?	             0@������������������������       �                     @�       �                   �^@8�Z$���?             *@������������������������       �                     @�       �                   Hp@����X�?             @������������������������       �                     @������������������������       �                      @�       �                    �?H�ՠ&��?             K@�       �                   �q@�t����?	             1@������������������������       �                     (@������������������������       �                     @�       �       	          ����?@-�_ .�?            �B@�       �                   �s@      �?
             0@�       �                   �a@��S�ۿ?	             .@������������������������       �                     &@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             5@�       �                    �?P����?             C@������������������������       �                     @�       �       	          033�?����X�?            �A@�       �                    �N@�����H�?	             2@������������������������       �                     &@�       �                    @O@����X�?             @������������������������       �                     �?�       �                    a@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �M@��.k���?	             1@������������������������       �                     @�       �                    �?ףp=
�?             $@�       �                     P@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       �z@     �~@     �X@     @z@      L@     �w@      6@      9@      @      4@      @       @              �?      @      �?      @              �?      �?              �?      �?               @      2@      �?      �?      �?                      �?      �?      1@      �?      @              @      �?                      (@      0@      @      0@      �?      (@              @      �?      @              �?      �?      �?                      �?              @      A@     0v@      (@     �B@              3@      (@      2@      (@      *@              @      (@      @      @              @      @      @      @      @              �?      @      �?       @               @      �?                      @              �?              @      6@     �s@      3@     �s@      �?              2@     �s@      &@     �V@      &@     �S@      @      O@      @      ?@      @      ?@       @      @       @       @       @                       @               @       @      ;@      �?              �?      ;@              .@      �?      (@      �?                      (@      �?                      ?@      @      1@      @      1@              $@      @      @      @       @      �?       @               @      �?               @                      @      @                      (@      @     �k@      @      ;@      @      $@      @      @              @      @                      @              1@      @     `h@       @      e@       @      O@              >@       @      @@              ,@       @      2@      �?              �?      2@      �?       @               @      �?                      0@             �Z@       @      :@              3@       @      @              @       @              @      @      @      �?              �?      @                      @      E@      D@      E@     �@@      @      0@      @       @      �?       @      �?                       @       @              �?      ,@              *@      �?      �?      �?                      �?      C@      1@      (@      0@      (@       @       @      �?      @              �?      �?              �?      �?              @      @      @      �?              �?      @              �?      @              @      �?                       @      :@      �?      6@              @      �?      @              �?      �?      �?                      �?              @     �t@     @Q@     p@      9@     `n@      (@      :@      @      �?      �?              �?      �?              9@      @      9@       @      @       @      @              �?       @               @      �?              5@                      �?      k@       @      @      @      @      �?      @                      �?              @     �j@      @     �h@      @     @X@              Y@      @     �I@             �H@      @               @     �H@       @      @      �?      @                      �?     �F@      �?      *@      �?      (@              �?      �?      �?                      �?      @@              1@              ,@      *@              "@      ,@      @      �?      @      �?                      @      *@             �R@      F@     �N@      3@      ,@      (@      @      @      @       @               @      @                      @      &@      @              @      &@       @      @              @       @      @                       @     �G@      @      (@      @      (@                      @     �A@       @      ,@       @      ,@      �?      &@              @      �?      @                      �?              �?      5@              *@      9@      @              $@      9@       @      0@              &@       @      @      �?              �?      @              @      �?               @      "@      @              �?      "@      �?      @              @      �?                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��^hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKᅔh~�B81         `       	          ����?�ڰ����?I           ��@       M                    �?������?!           0|@                          �c@0�����?�            �x@              
             �?b����o�?(            �R@������������������������       �                    �H@                           �?$��m��?             :@       
                    �?�<ݚ�?             "@       	                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @                          `c@�t����?
             1@������������������������       �        	             .@������������������������       �                      @       ,       
             �?��+Q���?�            0t@                           �?�d�K���?'            �P@              	          ����?�GN�z�?             6@                           ^@      �?             @������������������������       �                     �?������������������������       �                     @              	          833�?�����H�?             2@������������������������       �                     @                          �b@r�q��?             (@                           _@�C��2(�?             &@������������������������       �                     @                           `@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?                           �?�<ݚ�?            �F@������������������������       �                     7@        +                    �?�eP*L��?             6@!       *       	          @33�?j���� �?             1@"       )                   �e@      �?
             ,@#       $                   �n@�q�q�?	             (@������������������������       �                     @%       &                   �b@r�q��?             @������������������������       �                     @'       (                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @-       >                    @L@     ��?�             p@.       7                   �h@@	tbA@�?�            �i@/       0                   �c@@9G��?            �H@������������������������       �                     =@1       6                   �h@ףp=
�?             4@2       5                    �?�}�+r��?             3@3       4                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             1@������������������������       �                     �?8       =                    �?@=��?k            �c@9       :                   hq@@4և���?
             ,@������������������������       �                     $@;       <                   �r@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        a             b@?       L                     P@�����?"            �H@@       K                    �?�d�����?             C@A       B                   �a@�t����?             A@������������������������       �                     2@C       F                   �l@      �?             0@D       E                    b@����X�?             @������������������������       �                     @������������������������       �                      @G       J                   �^@�����H�?             "@H       I                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     &@N       U                    I@r�z-��?'            �J@O       T                    @N@      �?             0@P       S                   �]@؇���X�?             @Q       R       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@V       Y                   �b@��%��?            �B@W       X       
             �?�	j*D�?             :@������������������������       �                     2@������������������������       �                      @Z       [                   �h@"pc�
�?             &@������������������������       �                     �?\       _                   Pd@ףp=
�?             $@]       ^                    �J@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @a       �                    �?�f��9��?(           0}@b       �                    �?LGz���?y             h@c       �                   �b@XKu"�<�?R            �_@d       e       	             �?|��?���?&             K@������������������������       �                     @f                           �Q@��C���?             �G@g       r                   Pl@�q�q�?             E@h       q                    @R���Q�?             4@i       j                    `@�KM�]�?             3@������������������������       �                     (@k       l                   ``@����X�?             @������������������������       �                     �?m       n                    �?r�q��?             @������������������������       �                     @o       p       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?s       t                   �o@      �?             6@������������������������       �                     @u       x                    @K@b�2�tk�?             2@v       w                   �p@      �?              @������������������������       �                     @������������������������       �                     @y       ~                   �e@z�G�z�?             $@z       {                   @_@�����H�?             "@������������������������       �                     @|       }       	          ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	          `ff@v���a�?,            @R@�       �                    �?�qM�R��?&            �P@�       �                    �F@����X�?             ,@������������������������       �                     @�       �                   `d@      �?              @������������������������       �                     @�       �                   pe@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	          `ff�?�&=�w��?            �J@������������������������       �        	             0@�       �                    �L@@-�_ .�?            �B@�       �                   �d@�g�y��?             ?@������������������������       �                     3@�       �       
             �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�       �                    �?r�q��?             @�       �       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �f@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?r�q��?'            �P@�       �                   �w@�8��8��?             H@�       �                   �j@����?�?            �F@������������������������       �                    �B@�       �                    �?      �?              @�       �                   ``@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   �q@b�2�tk�?             2@�       �                    @J@8�Z$���?             *@������������������������       �                     @�       �                   �a@z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�u����?�             q@�       �                    �?`�q��־?�             m@�       �       	          ����?д>��C�?             =@������������������������       �                     @�       �                   `\@$�q-�?             :@�       �       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �J@�nkK�?             7@�       �                    �I@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@�       �       	          033�?@��j$޷?�            �i@�       �                   �k@�k~X��?/             R@������������������������       �                     B@�       �                   �l@������?             B@������������������������       �                     �?������������������������       �                    �A@�       �       
             �?t��ճC�?R            �`@�       �                   Pb@��7�K¨?L            @^@�       �                    �R@���1��?D            �Z@������������������������       �        B            �Y@�       �                   �b@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    \@؇���X�?             ,@������������������������       �                     �?�       �                    �?$�q-�?             *@�       �                    �F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�       �                   @_@�eP*L��?             &@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �       	              @���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �h@��]�T��?            �D@�       �                    �M@ףp=
�?	             $@������������������������       �                     @�       �                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �b@`՟�G��?             ?@�       �                   �[@`�Q��?             9@������������������������       �                     @�       �                    �?��s����?             5@������������������������       �                      @�       �       	          ����?�KM�]�?             3@������������������������       �                      @������������������������       �                     1@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B        {@     @~@     s@     @b@     �q@     �[@      1@      M@             �H@      1@      "@       @      @       @       @       @                       @              @      .@       @      .@                       @     �p@     �J@      ;@      D@      1@      @      �?      @      �?                      @      0@       @      @              $@       @      $@      �?      @              @      �?              �?      @                      �?      $@     �A@              7@      $@      (@      $@      @      @      @      @      @      @              �?      @              @      �?      �?      �?                      �?               @      @                      @     `n@      *@     �i@      @     �G@       @      =@              2@       @      2@      �?      �?      �?              �?      �?              1@                      �?     �c@      �?      *@      �?      $@              @      �?              �?      @              b@             �C@      $@      <@      $@      8@      $@      2@              @      $@      @       @      @                       @      �?       @      �?      �?      �?                      �?              @      @              &@              2@     �A@      �?      .@      �?      @      �?      �?              �?      �?                      @              "@      1@      4@       @      2@              2@       @              "@       @              �?      "@      �?      @      �?              �?      @              @              `@      u@     �X@     �W@      V@     �C@      :@      <@      @              3@      <@      ,@      <@      @      1@       @      1@              (@       @      @      �?              �?      @              @      �?      �?      �?                      �?      �?              &@      &@      @              @      &@      @      @              @      @               @       @      �?       @              @      �?      @      �?                      @      �?              @              O@      &@     �N@      @      $@      @      @              @      @      @              �?      @              @      �?             �I@       @      0@             �A@       @      >@      �?      3@              &@      �?              �?      &@              @      �?      �?      �?      �?                      �?      @              �?      @              @      �?              &@     �K@      @      F@      �?      F@             �B@      �?      @      �?      @      �?                      @              @      @              @      &@       @      &@              @       @       @               @       @              @              >@     �n@      .@     @k@      @      8@      @               @      8@      �?       @      �?                       @      �?      6@      �?       @               @      �?                      ,@      $@     @h@      �?     �Q@              B@      �?     �A@      �?                     �A@      "@     �^@      @     �]@      �?     �Z@             �Y@      �?      @              @      �?               @      (@      �?              �?      (@      �?      �?              �?      �?                      &@      @      @      @              @      @              @      @       @      @                       @      .@      :@      �?      "@              @      �?       @               @      �?              ,@      1@       @      1@      @              @      1@       @               @      1@       @                      1@      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJB�PhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �                    �?�LT ���?N           ��@       O       	          033�?����:�?B           �~@       D                    �?p�ݯ��?�             j@              
             �?8�����?i            �b@                           �?D˩�m��?5            �R@                           �?0,Tg��?             E@                           �?      �?             @������������������������       �                      @	       
                   `_@      �?              @������������������������       �                     �?������������������������       �                     �?              	          ����?���y4F�?             C@������������������������       �                     >@������������������������       �                      @                          @e@     ��?             @@                           �F@ܷ��?��?             =@                           �E@�q�q�?             @������������������������       �                     �?                          �b@      �?              @������������������������       �                     �?������������������������       �                     �?                          �_@$�q-�?             :@������������������������       �                     "@                          �[@�t����?             1@                          �Y@����X�?             @������������������������       �                     @                           b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@������������������������       �                     @        /                   pc@���!pc�?4            @S@!       .       	          ����?��2(&�?             F@"       -                   �f@X�EQ]N�?            �E@#       &                    �?�����?             E@$       %                   `^@���Q��?             @������������������������       �                      @������������������������       �                     @'       (                    �?�?�|�?            �B@������������������������       �                     >@)       ,                   �a@؇���X�?             @*       +                   @b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?0       =                   Pd@�eP*L��?            �@@1       6                   `o@�q�q�?             2@2       3                   d@�����H�?             "@������������������������       �                     @4       5                   @_@      �?             @������������������������       �                     �?������������������������       �                     @7       <                    d@X�<ݚ�?             "@8       9                    �?r�q��?             @������������������������       �                     @:       ;                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @>       ?                    �L@z�G�z�?	             .@������������������������       �                      @@       C                    �?և���X�?             @A       B                   f@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @E       N       	          833�? 	��p�?#             M@F       G       
             �?���}<S�?             G@������������������������       �                     A@H       K                    �?�q�q�?             (@I       J                   ``@�q�q�?             @������������������������       �                     @������������������������       �                      @L       M                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     (@P       o       	          ����?�ӖF2��?�            �q@Q       R                   �Q@д>��C�?*             M@������������������������       �                      @S       d                    �?؇���X�?)             L@T       U       	          `ff�?@4և���?             E@������������������������       �                     @V       c                   �o@$�q-�?            �C@W       \                    �? �Cc}�?             <@X       Y                   @_@      �?             @������������������������       �                     �?Z       [                     L@�q�q�?             @������������������������       �                     �?������������������������       �                      @]       b                    �? �q�q�?             8@^       a                   �W@@4և���?
             ,@_       `                   �a@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@������������������������       �                     $@������������������������       �        	             &@e       f                   �Y@X�Cc�?
             ,@������������������������       �                     @g       l                   @^@X�<ݚ�?             "@h       k                   �[@      �?             @i       j       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @m       n                    �H@z�G�z�?             @������������������������       �                     �?������������������������       �                     @p       }                    _@ \sF��?�            @l@q       z                   �^@ܷ��?��?"             M@r       s                    _@�>����?              K@������������������������       �                     9@t       y                   �j@\-��p�?             =@u       x                     K@���|���?	             &@v       w                   �g@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@{       |                    �J@      �?             @������������������������       �                      @������������������������       �                      @~       �                    `R@�Ń��̧?j             e@       �                    @M@ ���+�?h            �d@������������������������       �        =             X@�       �       	          ����?hA� �?+            �Q@�       �                   xu@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    c@Pa�	�?'            �P@�       �       	          033�?0�)AU��?             �L@������������������������       �                     8@�       �                    �?Pa�	�?            �@@������������������������       �                     &@�       �                    �M@���7�?             6@������������������������       �                     �?������������������������       �                     5@�       �                   �`@�����H�?             "@�       �                   �c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?��De�h�?           �z@�       �                    @L@kI.!��?�            `u@�       �                    @ĴF���?�            �n@�       �                   @c@�8��!�?�             l@�       �                    �?և���X�?	             ,@������������������������       �                     @�       �                   �K@���Q��?             $@������������������������       �                     @�       �                   �\@և���X�?             @������������������������       �                     @�       �                   `X@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   pk@h+�"��?�            `j@�       �       	          ����?�L��ȕ?;            @W@������������������������       �        :             W@������������������������       �                     �?�       �       
             �?�1e�3��?F            �]@�       �                    ]@�+e�X�?             9@�       �                   pf@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?ףp=
�?             4@�       �                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     1@�       �                   @[@�L��ȕ?5            @W@�       �                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        3            �V@�       �                   �c@�q�q�?             5@������������������������       �                     @�       �                   �`@@�0�!��?             1@������������������������       �                     �?�       �                    �F@      �?
             0@�       �       
             �?      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    @O@�q�q�?@             X@�       �       	          ����?�p����?*            �N@�       �                   0a@�Gi����?            �B@�       �                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�       �       	          033�?� �	��?             9@�       �                    c@���|���?             6@�       �                    �L@X�<ݚ�?             2@�       �                   �a@      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?�z�G��?	             $@�       �                    @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    b@�q�q�?             8@������������������������       �                     $@�       �                    �?X�Cc�?
             ,@�       �                    @      �?              @������������������������       �                     @������������������������       �                     �?�       �       	          ���@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �       
             �?b�h�d.�?            �A@�       �       	          ����?�eP*L��?             &@������������������������       �                     @�       �       	          033@      �?              @������������������������       �                     @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �? �q�q�?             8@������������������������       �        
             4@�       �                    �?      �?             @������������������������       �                      @�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?�             
             �?F~��7�?4            �T@�       �                   �n@���!pc�?(            �P@�       �                    �?H�z�G�?             D@������������������������       �                     @�       �                    �?�!���?             A@�       �       	          @33�?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �N@d}h���?             <@�       �                   �`@�q�q�?             2@������������������������       �                      @�       �                   �[@���Q��?             $@������������������������       �                      @�       �                    @      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     $@�                          �? ��WV�?             :@�       �                    �?      �?             0@������������������������       �                     @�       �                   �s@�C��2(�?             &@������������������������       �                      @�                          @[@�q�q�?             @������������������������       �                     �?            	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     1@�t�b��(     h�h(h+K ��h-��R�(KMKK��h_�BP       �y@     �@     @X@     �x@     @S@     �`@     @R@     �S@      1@     �L@      &@      ?@      @      �?       @              �?      �?              �?      �?               @      >@              >@       @              @      :@      @      :@      �?       @              �?      �?      �?              �?      �?               @      8@              "@       @      .@       @      @              @       @      �?       @                      �?              $@      @              L@      5@      C@      @      C@      @      C@      @       @      @       @                      @      B@      �?      >@              @      �?       @      �?              �?       @              @                      �?              �?      2@      .@      @      (@      �?       @              @      �?      @      �?                      @      @      @      @      �?      @              �?      �?              �?      �?                      @      (@      @       @              @      @       @      @              @       @               @              @      K@      @      E@              A@      @       @       @      @              @       @               @      @       @                      @              (@      4@     �p@      $@      H@       @               @      H@      @     �C@              @      @      B@      @      9@       @       @      �?              �?       @      �?                       @      �?      7@      �?      *@      �?      @              @      �?                      $@              $@              &@      @      "@              @      @      @      �?      @      �?      �?      �?                      �?               @      @      �?              �?      @              $@      k@      @      J@      @      I@              9@      @      9@      @      @      �?      @              @      �?              @                      2@       @       @       @                       @      @     �d@      @     `d@              X@      @     �P@      �?      @              @      �?               @      P@      �?      L@              8@      �?      @@              &@      �?      5@      �?                      5@      �?       @      �?      @      �?                      @              @      �?      �?              �?      �?             �s@     @[@     �q@     �N@      l@      5@     `j@      ,@       @      @      @              @      @              @      @      @      @              �?      @      �?                      @     `i@       @      W@      �?      W@                      �?     �[@      @      3@      @      �?      @              @      �?              2@       @      �?       @               @      �?              1@              W@      �?      �?      �?      �?                      �?     �V@              ,@      @              @      ,@      @              �?      ,@       @      @       @               @      @               @              L@      D@      ;@      A@      6@      .@      &@      �?      &@                      �?      &@      ,@       @      ,@       @      $@      �?      @              @      �?              @      @      @       @      @                       @              �?              @      @              @      3@              $@      @      "@      �?      @              @      �?              @       @      @                       @      =@      @      @      @              @      @       @      @              �?       @      �?                       @      7@      �?      4@              @      �?       @              �?      �?              �?      �?             �A@      H@      2@      H@      1@      7@      @              &@      7@      @      �?              �?      @              @      6@      @      (@               @      @      @       @              @      @      @                      @              $@      �?      9@      �?      .@              @      �?      $@               @      �?       @              �?      �?      �?      �?                      �?              $@      1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ;�}hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �                    �?��+�?J           ��@       9       	          ����?rn�#���?<            @       4                    �?V1���?r             e@              
             �?d�
��?Y            �`@                          �`@Ԫ2��?&            �L@              	          ����?x�����?            �C@������������������������       �                     :@                          `_@�n_Y�K�?             *@	                           �O@      �?              @
                          �Z@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     2@       )                    �L@������?3            �R@       &       	             �?f1r��g�?&            �J@                          pc@H%u��?#             I@������������������������       �                     >@       #                    �?�z�G��?             4@                            �I@�E��ӭ�?             2@                           �?z�G�z�?             .@                          �c@����X�?             @������������������������       �                     �?                          �f@r�q��?             @                           e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                          pf@      �?              @������������������������       �                     @������������������������       �                     �?!       "                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?$       %                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?'       (                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?*       3                    �?�eP*L��?             6@+       0                    �?�q�q�?
             2@,       /                     P@      �?             $@-       .                   �`@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @1       2                   �p@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @5       8                    �?�?�|�?            �B@6       7       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     >@:       I                    �?��=���?�            �t@;       B                   xr@�z�G��?             D@<       A                    �J@�J�4�?             9@=       >       
             �?�q�q�?             @������������������������       �                      @?       @                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     3@C       H                   pc@��S���?             .@D       E                   s@���|���?             &@������������������������       �                     @F       G                   `\@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @J       }                   �z@��m���?�            r@K       |       	          `ff@ �媩��?�            �q@L       Q                    Z@ �q�q�?�            �p@M       N                   Pd@z�G�z�?             $@������������������������       �                     @O       P                   a@�q�q�?             @������������������������       �                     �?������������������������       �                      @R       {       	          `ff @�)���?�            �o@S       Z                   �[@0z�(>��?�            �j@T       U                     J@�����?             5@������������������������       �                     "@V       Y                    �?r�q��?             (@W       X                   �k@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @[       r                   0c@�q�q��?t             h@\       o                    �R@��$����?i            �e@]       n                   ``@`��>�ϗ?g            @e@^       m                    �?      �?(             P@_       l       
             �?@9G��?            �H@`       i                   Xr@`Ӹ����?            �F@a       h       	          ����? qP��B�?            �E@b       g                   l@�8��8��?             (@c       d                    �?r�q��?             @������������������������       �                     @e       f                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     ?@j       k                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     .@������������������������       �        ?            �Z@p       q                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?s       t                   `c@z�G�z�?             4@������������������������       �                     @u       v       	          033�?�IєX�?	             1@������������������������       �                     "@w       x                   pl@      �?              @������������������������       �                     @y       z                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                    �D@������������������������       �                     5@~                          �_@      �?             @������������������������       �                      @������������������������       �                      @�       �       
             �?8	C)��?           @z@�       �                   a@����"�?n            �e@�       �                    �?��oh���?0            @R@�       �                   �r@���@M^�?             ?@�       �                    �?J�8���?             =@�       �                   `Z@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    @L@"pc�
�?             6@�       �                   pb@�q�q�?             "@�       �                    @K@      �?              @�       �                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �^@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    `@$�q-�?
             *@������������������������       �                     &@�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    \@�����?             E@�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �s@@-�_ .�?            �B@������������������������       �                    �@@�       �                   @[@      �?             @������������������������       �                     �?�       �                    �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @K@��j2��?>            @Y@�       �                    �?:���W�?$            �M@������������������������       �                     ,@�       �                    �?��S���?            �F@�       �                    @v�2t5�?            �D@�       �                   �`@^H���+�?            �B@�       �                    �G@      �?             <@�       �                    �?      �?
             0@�       �       	              @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@�       �                   �d@      �?             (@�       �                   �\@      �?              @������������������������       �                     @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �I@�q�q�?             "@�       �                   `a@؇���X�?             @�       �                    d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?����X�?             E@�       �                   �_@�q�q�?             (@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   Pr@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   Pa@�������?             >@������������������������       �                      @�       �       
             �?�>4և��?             <@������������������������       �                     �?�       �                    �?PN��T'�?             ;@�       �       	          `ff�?�C��2(�?             6@�       �                   �k@؇���X�?             ,@������������������������       �                     $@�       �                   �l@      �?             @������������������������       �                     �?�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    @���Q��?             @�       �       	          ����?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    @L@@;�"�?�            �n@�       �                    �?����?�            @i@������������������������       �        M            �^@�       �                   �_@86��Z�?5            �S@�       �                     I@�<ݚ�?             2@�       �                    @H@      �?              @�       �                    Y@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     $@�       �       	          ����?��v$���?*            �N@�       �                    @G@ qP��B�?            �E@������������������������       �                     6@�       �                    �G@���N8�?             5@�       �                    �?z�G�z�?             @������������������������       �                     @�       �                   @[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@������������������������       �                     2@�       �                    �?      �?             F@�       �                    �M@�����?             5@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                     R@�X�<ݺ?             2@������������������������       �                     ,@�       �                    `R@      �?             @������������������������       �                     �?������������������������       �                     @�             	          ����?�û��|�?             7@�                         ps@      �?             0@�                          �L@��S�ۿ?             .@             	          pff�?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             &@������������������������       �                     �?������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�BP       x@     ��@     @V@     �y@      P@     @Z@     �O@     @Q@       @     �H@       @      ?@              :@       @      @      @      @      �?      @      �?                      @       @              @                      2@     �K@      4@     �F@       @      F@      @      >@              ,@      @      *@      @      (@      @      @       @              �?      @      �?       @      �?       @                      �?      @              @      �?      @                      �?      �?       @               @      �?              �?      �?              �?      �?              �?       @               @      �?              $@      (@      @      (@      @      @      @      @              @      @               @              �?      @              @      �?              @              �?      B@      �?      @              @      �?                      >@      9@      s@      (@      <@      @      5@      @       @       @               @       @       @                       @              3@       @      @      @      @      @              �?      @      �?                      @      @              *@     @q@      &@      q@      &@     �o@       @       @              @       @      �?              �?       @              "@     �n@      "@     �i@       @      3@              "@       @      $@       @       @       @                       @               @      @      g@      @      e@       @      e@       @      O@       @     �G@       @     �E@      �?      E@      �?      &@      �?      @              @      �?       @      �?                       @              @              ?@      �?      �?      �?                      �?              @              .@             �Z@      �?      �?              �?      �?              @      0@      @              �?      0@              "@      �?      @              @      �?      �?      �?                      �?             �D@              5@       @       @               @       @             �r@      _@     �P@      [@      0@     �L@      (@      3@      $@      3@      @      �?              �?      @              @      2@      @      @      @      @      �?       @               @      �?               @      @       @                      @              �?      �?      (@              &@      �?      �?      �?                      �?       @              @      C@       @      @       @                      @       @     �A@             �@@       @       @              �?       @      �?              �?       @              I@     �I@      C@      5@      ,@              8@      5@      8@      1@      8@      *@      5@      @      .@      �?      �?      �?      �?                      �?      ,@              @      @      @       @      @               @       @       @                       @              @      @      @      �?      @      �?      �?      �?                      �?              @       @                      @              @      (@      >@      @      @      @       @               @      @              �?      @              @      �?              @      7@       @              @      7@      �?              @      7@       @      4@       @      (@              $@       @       @      �?              �?       @               @      �?                       @       @      @      �?      @      �?      �?      �?                      �?               @      �?             �l@      0@     �h@      @     �^@             �R@      @      ,@      @      @      @      @      �?              �?      @                      @      $@              N@      �?      E@      �?      6@              4@      �?      @      �?      @              �?      �?              �?      �?              0@              2@             �@@      &@      3@       @       @      �?       @                      �?      1@      �?      ,@              @      �?              �?      @              ,@      "@      ,@       @      ,@      �?      @      �?              �?      @              &@                      �?              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJw��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�:         b                   P`@2���xA�?:           ��@       3                    �?��$4d�?           �z@       &       
             �?��
ц��?k             e@                           �?&<k����?8            @V@       
                    �?�q�q�?             (@       	                    �?      �?              @              	          ����?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       #                    �Q@�s�c���?1            @S@              
             �?�ӖF2��?.            �Q@                           �M@���Q��?             @                           @I@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @                          �_@���7�?*            �P@                           �?@3����?"             K@������������������������       �                    �G@                           @؇���X�?             @                          `Z@z�G�z�?             @                           \@�q�q�?             @������������������������       �                     �?                          �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @               	             �?r�q��?             (@������������������������       �                     @!       "       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     @$       %                    �?      �?             @������������������������       �                     @������������������������       �                     @'       ,       	          ����?R���Q�?3             T@(       )                    �?��S�ۿ?)             N@������������������������       �        $             J@*       +                   @V@      �?              @������������������������       �                     @������������������������       �                     @-       .                    �?�z�G��?
             4@������������������������       �                     @/       0                   @d@@�0�!��?	             1@������������������������       �                     (@1       2       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @4       _       
             �?�}�}CS�?�            0p@5       V                   `_@ ,��-�?�            �m@6       E                   `Z@ؗp�'ʸ?x            �h@7       D                   �`@���c���?              J@8       =                   �_@R�}e�.�?             :@9       <                    \@�KM�]�?             3@:       ;       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@>       ?                    `@����X�?             @������������������������       �                     @@       A       	             �?      �?             @������������������������       �                     �?B       C                   l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     :@F       U       	          ����?@��8��?X             b@G       H                     K@�˹�m��?             C@������������������������       �                     .@I       T                    �?�LQ�1	�?             7@J       M                   �[@@�0�!��?             1@K       L                    �?      �?              @������������������������       �                     �?������������������������       �                     �?N       O                    �?�r����?             .@������������������������       �                     "@P       Q                   �\@�q�q�?             @������������������������       �                     �?R       S                   �c@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �        =            �Z@W       \                   `b@R���Q�?             D@X       Y                    @L@      �?             @@������������������������       �        
             4@Z       [                    �L@r�q��?             (@������������������������       �                      @������������������������       �                     $@]       ^                     I@      �?              @������������������������       �                     @������������������������       �                     @`       a       	            �?�û��|�?             7@������������������������       �                     "@������������������������       �        	             ,@c       �       	          033�?�::C��?3           �~@d       �                    �?��i,��?�            `x@e       |       
             �?���5��?\             a@f       g       	          ����?��$�4��?+            �M@������������������������       �                     4@h       i                   �`@�q�q�?            �C@������������������������       �                     @j       {                    �?�E��ӭ�?             B@k       x                    �?\X��t�?             7@l       o                   pb@���Q��?             4@m       n       	          033�?�����H�?             "@������������������������       �                      @������������������������       �                     �?p       q                    @D@���|���?             &@������������������������       �                     �?r       w                   �r@�z�G��?             $@s       v                    �?      �?             @t       u       	          hff�?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @y       z                    �K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@}       �                    �?v��:ө�?1            �S@~       �                   �f@l��
I��?             ;@       �                   Xv@�q�q�?             8@�       �                   �c@��2(&�?             6@������������������������       �                     *@�       �                    �?�q�q�?             "@�       �                   d@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?�\�u��?"            �I@�       �                   �Y@�<ݚ�?            �F@������������������������       �                     @�       �       	          ����?r�q��?             E@�       �                   ``@�p ��?            �D@�       �       	          ����?�����?             3@�       �                    �?     ��?             0@�       �       	          @33�?$�q-�?
             *@�       �                   @c@      �?              @������������������������       �                     @�       �                   d@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@������������������������       �                     �?������������������������       �                     @�       �       
             �?������?�            �o@�       �                    �?     ��?)             P@�       �                    �K@���y4F�?             3@������������������������       �        
             (@�       �                   �q@և���X�?             @�       �                   @a@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �_@�q�q�?            �F@�       �                    @և���X�?             5@�       �                    �A@�q�q�?
             2@������������������������       �                      @�       �       	          ����?      �?	             0@������������������������       �                     �?�       �                    �?z�G�z�?             .@�       �                   `c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          ����?�8��8��?             (@������������������������       �                     $@�       �                   m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �a@      �?             8@�       �                   �`@�q�q�?             @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �Z@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    @N@�X�<ݺ?	             2@������������������������       �                     &@�       �                    @؇���X�?             @������������������������       �                     @�       �                   �d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �d@�J�-/��?t            �g@�       �                   �s@�>����?G             [@�       �       	            �?P���Q�?B             Y@�       �                    �?�(\����?5             T@�       �                   �m@�����H�?             "@�       �                   pd@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   n@ ��PUp�?.            �Q@������������������������       �                     D@�       �       	          ����?�g�y��?             ?@�       �                    @F@XB���?             =@������������������������       �        	             1@�       �                    �?�8��8��?             (@������������������������       �                     $@�       �                   @Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   pa@R���Q�?             4@������������������������       �                     @�       �                    @�θ�?	             *@�       �       	          ����?r�q��?             (@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     �?�       �                    @L@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �        -            @T@�       �                    \@�\m����?:             Y@�       �                    �G@���Q��?             $@������������������������       �                      @�       �                   @[@      �?              @������������������������       �                     @�       �                   �a@���Q��?             @������������������������       �                      @������������������������       �                     @�                         g@ ��~���?4            �V@�       �                    _@      �?3             V@�       �                   �^@      �?             8@�       �       	          033@"pc�
�?             6@�       �       
             �?X�<ݚ�?             "@������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                      @�                          �M@     p�?'             P@�                          @��hJ,�?             A@�                          c@      �?             @@�       �                    �? �q�q�?             8@������������������������       �                     3@�                           �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @                         a@      �?              @                        Pm@z�G�z�?             @������������������������       �                     @������������������������       �                     �?                        �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?	      
                    K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     >@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KMKK��h_�B�       Px@     ��@     �Y@     Pt@     �S@     �V@      0@     @R@       @      @      @      @      @      �?      @                      �?              @      @               @     @Q@      @     �P@       @      @       @      �?              �?       @                       @      @     �O@      �?     �J@             �G@      �?      @      �?      @      �?       @              �?      �?      �?      �?                      �?               @               @       @      $@              @       @      @       @                      @      @      @              @      @              O@      2@      L@      @      J@              @      @              @      @              @      ,@      @              @      ,@              (@      @       @      @                       @      9@     @m@      0@     �k@      $@     @g@      @     �F@      @      3@       @      1@       @      �?              �?       @                      0@      @       @      @               @       @              �?       @      �?       @                      �?              :@      @     �a@      @     �A@              .@      @      4@      @      ,@      �?      �?      �?                      �?       @      *@              "@       @      @              �?       @      @              @       @                      @             �Z@      @      A@       @      >@              4@       @      $@       @                      $@      @      @      @                      @      "@      ,@      "@                      ,@     �q@     �i@     �p@     �^@      L@     @T@      *@      G@              4@      *@      :@      @              $@      :@      $@      *@       @      (@      �?       @               @      �?              @      @              �?      @      @      @      @       @      @       @                      @      �?              @               @      �?       @                      �?              *@     �E@     �A@       @      3@      @      3@      @      3@              *@      @      @      @      @      @                      @              @       @              @             �A@      0@     �A@      $@              @     �A@      @     �A@      @      *@      @      *@      @      (@      �?      @      �?      @              @      �?              �?      @              @              �?       @               @      �?                      @      6@                      �?              @     `j@      E@      >@      A@      .@      @      (@              @      @      �?      @              @      �?               @              .@      >@      (@      "@      (@      @               @      (@      @              �?      (@      @      �?       @      �?                       @      &@      �?      $@              �?      �?      �?                      �?              @      @      5@       @      @      �?      �?              �?      �?              �?      @      �?                      @      �?      1@              &@      �?      @              @      �?       @      �?                       @     �f@       @      Y@       @     �W@      @     �S@       @       @      �?       @      �?       @                      �?      @             �Q@      �?      D@              >@      �?      <@      �?      1@              &@      �?      $@              �?      �?      �?                      �?       @              1@      @      @              $@      @      $@       @       @       @               @       @               @                      �?      @      @      @                      @     @T@              3@     @T@      @      @               @      @       @      @              @       @               @      @              *@     @S@      &@     @S@      @      2@      @      2@      @      @              @      @      �?      @                      �?              *@       @              @     �M@      @      =@      @      <@      �?      7@              3@      �?      @      �?                      @      @      @      �?      @              @      �?               @      �?       @                      �?      �?      �?              �?      �?                      >@       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ[��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�8         �                    �?��IT�?J           ��@       �                    �?t>UhVJ�?C           p@       P                    �?r٣����?�            �v@                           �?�8p/�5�?`            �a@                          �f@:�&���?            �C@              	            �?$G$n��?            �B@                          d@     ��?             0@                          �c@      �?	             $@	                          �r@����X�?             @
                          �[@r�q��?             @                          g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     5@������������������������       �                      @       O                   �w@h0�����?G            @Y@                           �?r�q��?D             X@              	          `ff�?$�q-�?
             *@                           �B@؇���X�?             @������������������������       �                     @                           Z@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       D                    �?��q7L��?:            �T@       A       	          ����?\X��t�?0            @Q@       ,                   ``@      �?)             M@        %                     J@"pc�
�?             6@!       $                   ``@      �?             @"       #                    �G@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @&       '                   �`@      �?             0@������������������������       �                     "@(       +                   0a@؇���X�?             @)       *                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @-       :                    e@<ݚ)�?             B@.       5                   �_@d}h���?             <@/       0                    a@�t����?             1@������������������������       �                     @1       4                   �^@�n_Y�K�?	             *@2       3       
             �?���!pc�?             &@������������������������       �                     @������������������������       �                      @������������������������       �                      @6       9       
             �?�C��2(�?             &@7       8                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @;       <                    �D@      �?              @������������������������       �                     @=       @                   �`@      �?             @>       ?                     G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @B       C       
             �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?E       N                   h@����X�?
             ,@F       G       
             �?և���X�?             @������������������������       �                     �?H       M                   �U@�q�q�?             @I       J                   `Y@      �?             @������������������������       �                     �?K       L       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @Q       v       	          ����?���K��?�            �k@R       [                    @K@@�҇��?5            �W@S       V                    �?X�EQ]N�?            �E@T       U                   �p@      �?              @������������������������       �                     @������������������������       �                     @W       X                   �a@ >�֕�?            �A@������������������������       �                     ?@Y       Z                   �n@      �?             @������������������������       �                      @������������������������       �                      @\       e                   @i@ҳ�wY;�?             �I@]       d       	             �?HP�s��?             9@^       _                   �[@�r����?             .@������������������������       �                     $@`       a       
             �?���Q��?             @������������������������       �                     �?b       c                    V@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        	             $@f       u                     P@�n_Y�K�?             :@g       h                    �?���N8�?             5@������������������������       �                     @i       p       
             �?�����H�?	             2@j       k                   �`@$�q-�?             *@������������������������       �                     $@l       o                    d@�q�q�?             @m       n                     L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?q       r                   �r@z�G�z�?             @������������������������       �                     @s       t                   �s@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @w       �                   �i@ �#�Ѵ�?U             `@x       y                    �?$G$n��?            �B@������������������������       �                     �?z              	          ����?�����H�?             B@{       ~       
             �?և���X�?             @|       }                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     =@�       �       	          033@�����?;             W@������������������������       �        /            @S@�       �                     K@��S�ۿ?             .@�       �       	             @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �                    �R@h�����?Y            �a@�       �                    �?��*����?X            `a@�       �       	          ����?"pc�
�?             6@�       �                    Z@�	j*D�?             *@������������������������       �                     @�       �       	          433�?ףp=
�?             $@�       �                   m@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@������������������������       �        I            @]@������������������������       �                     �?�       �                    `@��B�}M�?           �y@�       �                    �?���
��??            �Z@�       �                   @c@,�|%�v�?2            @U@�       �                    `Q@�>4և��?             <@�       �                    �?�8��8��?             8@�       �                   @_@z�G�z�?             $@������������������������       �                     @�       �                   0a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �        	             ,@�       �                    �R@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �L@P̏����?!            �L@������������������������       �                     :@�       �                    �?`՟�G��?             ?@������������������������       �                     (@�       �                    �P@�d�����?             3@�       �                    �?�n_Y�K�?
             *@�       �                    �?z�G�z�?             @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �r@      �?              @������������������������       �                     @�       �                   @[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?���7�?             6@������������������������       �                     (@�       �                   �o@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �       
             �?�GN�z�?�            @s@�       �                    �?�~8�e�?@            �Y@�       �       	             �?��X��?             <@�       �                     G@�G�z��?             4@������������������������       �                     $@�       �                   hq@ףp=
�?             $@�       �                    �N@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?~�hP��?0            �R@�       �                    �?\X��t�?             7@�       �                   �p@D�n�3�?             3@�       �                    �K@ҳ�wY;�?             1@������������������������       �                     @�       �                    @���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   Pn@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?������?            �I@�       �       	          `ff�?V������?            �B@�       �                   `]@�\��N��?             3@�       �       	          @33�?؇���X�?             @������������������������       �                     @�       �                   @Z@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          ����?�q�q�?             (@������������������������       �                      @�       �                    �I@z�G�z�?             $@�       �                    �F@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�����H�?             2@�       �       	             
@r�q��?             (@�       �                   �^@ףp=
�?             $@������������������������       �                     @�       �                   �k@      �?             @������������������������       �                      @�       �                    @M@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   @e@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?�       �                    �L@p�eU}�?�            �i@�       �                   �O@@]����?t            @f@�       �                    �F@      �?              @������������������������       �                     @�       �                    �J@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   @g@`��>�ϗ?q            @e@������������������������       �        p             e@������������������������       �                      @�              	          ����?      �?             <@�       �                    @M@�����?             5@�       �                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @t@�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?                         �?����X�?             @������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�B0       �w@     Ѐ@     @W@     �y@      V@     0q@     �M@     @T@      @      @@      @      @@      @      &@      @      @       @      @      �?      @      �?      �?              �?      �?                      @      �?              @                      @              5@       @              J@     �H@      J@      F@      (@      �?      @      �?      @              @      �?              �?      @              @              D@     �E@      >@     �C@      =@      =@      @      2@      @      @      @      �?              �?      @                       @      �?      .@              "@      �?      @      �?      �?      �?                      �?              @      9@      &@      6@      @      (@      @      @               @      @       @      @              @       @                       @      $@      �?       @      �?       @                      �?       @              @      @              @      @      �?      �?      �?      �?                      �?       @              �?      $@              $@      �?              $@      @      @      @      �?               @      @       @       @              �?       @      �?              �?       @                       @      @                      @      =@     @h@      7@     �Q@      @      C@      @      @      @                      @       @     �@@              ?@       @       @       @                       @      2@     �@@       @      7@       @      *@              $@       @      @              �?       @       @       @                       @              $@      0@      $@      0@      @              @      0@       @      (@      �?      $@               @      �?      �?      �?      �?                      �?      �?              @      �?      @              �?      �?              �?      �?                      @      @     �^@      @      @@      �?              @      @@      @      @       @      @              @       @               @                      =@      �?     �V@             @S@      �?      ,@      �?      @      �?                      @              $@      @     �`@      @     �`@      @      2@      @      "@      @              �?      "@      �?      @      �?                      @              @              "@             @]@      �?             �q@      `@     �H@      M@      H@     �B@      @      7@       @      6@       @       @              @       @       @       @                       @              ,@      @      �?      @                      �?     �E@      ,@      :@              1@      ,@      (@              @      ,@      @       @      @      �?      �?      �?      �?                      �?      @              �?      @              @      �?      �?              �?      �?                      @      �?      5@              (@      �?      "@              "@      �?             �m@     �Q@      F@      M@      3@      "@      &@      "@      $@              �?      "@      �?      @              @      �?                      @       @              9@     �H@      *@      $@      &@       @      &@      @      @              @      @              @      @                       @       @       @       @                       @      (@     �C@      &@      :@      "@      $@      �?      @              @      �?       @      �?                       @       @      @               @       @       @       @       @       @                       @      @               @      0@       @      $@      �?      "@              @      �?      @               @      �?      �?      �?                      �?      �?      �?      �?                      �?              @      �?      *@              *@      �?             @h@      (@     �e@      @      @      @      @               @      @              @       @              e@       @      e@                       @      5@      @      3@       @       @      �?              �?       @              1@      �?      1@                      �?       @      @       @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�m]hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B6         �       
             �?��IT�?B           ��@       W                    �?H�,�7��?X           8�@                           �?�}��?�            �m@              	          ���@�w��#��?             I@                          `X@���j��?             G@������������������������       �                     @                          �Q@>��C��?            �E@������������������������       �                     @	                          @q@z�G�z�?             D@
                           �?�t����?             A@              	          ����?      �?             @@������������������������       �        	             .@                          `c@�t����?             1@                           b@      �?
             0@������������������������       �                     *@              
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                           @L@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @       *                   P`@��3E��?u            @g@                           �?x�G�z�?3             T@                           �?����e��?)            �P@������������������������       �        !            �L@              
             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @        )                    @؇���X�?
             ,@!       (                   @L@�<ݚ�?             "@"       #                    \@�q�q�?             @������������������������       �                     �?$       %                   �^@���Q��?             @������������������������       �                     �?&       '                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @+       T                   �f@�e�}|�?B            �Z@,       7                    �?zP1�??            @Y@-       0                   �^@�8��8��?             B@.       /                    a@r�q��?
             (@������������������������       �                      @������������������������       �        	             $@1       6                    �? �q�q�?             8@2       5       	          ����?�����H�?             "@3       4                    �J@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@8       9       
             �?�7�֥��?'            @P@������������������������       �                     @:       M                   ``@ 1_#�?#            �M@;       <                   �a@j���� �?             A@������������������������       �                      @=       H                    `@��
ц��?             :@>       G       	          ���@b�2�tk�?             2@?       F                   (q@��
ц��?             *@@       E                   pc@���|���?             &@A       D                    _@և���X�?             @B       C                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @I       L                    �?      �?              @J       K                   0b@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @N       O                   Pa@�J�4�?             9@������������������������       �                     @P       Q                    d@���7�?             6@������������������������       �        
             3@R       S       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?U       V       	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @X       m                    @G@|fG�b�?�            �s@Y       f                   Pb@��d��?'            �O@Z       [                   �_@��S�ۿ?            �F@������������������������       �                     3@\       e                    �?ȵHPS!�?             :@]       `                    `@     ��?
             0@^       _                    �C@�q�q�?             @������������������������       �                     �?������������������������       �                      @a       b                   �l@$�q-�?             *@������������������������       �                     "@c       d                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@g       h                    �?b�2�tk�?
             2@������������������������       �                     @i       l                   �l@�8��8��?             (@j       k                   �j@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@n       �                   `_@$Q�q�?�            �o@o       p                    @K@�Q��k�?b             d@������������������������       �                    �H@q       �       	          ����?�g+��@�?E            �[@r       �                   �a@���c���?             J@s       t       	          ����?��G���?            �B@������������������������       �                     *@u       v                    �K@�q�q�?             8@������������������������       �                      @w       ~                    �O@�GN�z�?             6@x       }                    @N@؇���X�?
             ,@y       |                   �`@"pc�
�?             &@z       {                    e@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @       �                    �?      �?              @�       �                    `@����X�?             @�       �                    _@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �        
             .@������������������������       �        &            �M@�       �                   �_@�ܸb���?;             W@�       �                   �^@�q�q�?             @������������������������       �                     �?�       �                    @L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?����"$�?6            �U@�       �                    @H@���5��?&            �L@������������������������       �                     �?�       �                   �`@ �Cc}�?%             L@������������������������       �        	             0@�       �                    �J@R���Q�?             D@�       �                    l@      �?              @�       �       	          `ff@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @     ��?             @@�       �                    �?(;L]n�?             >@������������������������       �                     :@�       �                   pa@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     =@�       �                    �?�Z{����?�            �v@�       �       	          ����?~��l��?O            �\@�       �                    �?� �	��?E             Y@�       �                    P@���=A�?3             S@�       �                    @O@     ��?	             0@�       �                    �?@4և���?             ,@�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                      @�       �                   �k@z�G�z�?*             N@�       �                    �?�}�+r��?             3@�       �                    �?      �?             @�       �                    ]@�q�q�?             @�       �                   Pa@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     .@�       �                   �b@���� �?            �D@�       �                    �?�}�+r��?             3@�       �                   pa@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             0@�       �                    �L@�eP*L��?             6@�       �                    ]@�q�q�?             2@�       �                   �[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   pf@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @������������������������       �                     @�       �                   �s@�q�q�?             8@�       �                   Pk@ףp=
�?             4@�       �                    �?8�Z$���?
             *@�       �                   �d@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �J@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �e@z�G�z�?
             .@�       �                    @N@$�q-�?	             *@�       �                   �a@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �       	             @�����?�            �o@�       �                    I@$�q-�?�            �n@�       �                    �N@�n_Y�K�?             *@������������������������       �                     @�       �       	          ����?      �?             $@�       �                   �b@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �_@0��d��?�            @m@�       �                   @c@     ��?             @@������������������������       �                     @�       �                    �L@ܷ��?��?             =@������������������������       �                     8@�       �                    q@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   xt@����?            @i@�       �                   �g@����e��?|            �h@�       �                    @L@@uvI��?z            �h@������������������������       �        f            `d@�       �                    �L@�FVQ&�?            �@@������������������������       �                      @������������������������       �                     ?@�       �                    �D@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�t�b�v     h�h(h+K ��h-��R�(KK�KK��h_�Bp       �w@     Ѐ@     @W@     �|@     �P@      e@     �@@      1@     �@@      *@              @     �@@      $@              @     �@@      @      >@      @      >@       @      .@              .@       @      .@      �?      *@               @      �?       @                      �?              �?               @      @      @              @      @                      @      A@      c@      @     @S@      �?     @P@             �L@      �?       @      �?                       @       @      (@       @      @       @      @              �?       @      @      �?              �?      @      �?                      @              @              @      ?@     �R@      ;@     �R@      @     �@@       @      $@       @                      $@      �?      7@      �?       @      �?      @              @      �?                      @              .@      8@     �D@      @              2@     �D@      ,@      4@               @      ,@      (@      @      &@      @      @      @      @      @      @      @      �?      @                      �?              @      @                       @              @      @      �?      @      �?              �?      @              @              @      5@      @              �?      5@              3@      �?       @               @      �?              @      �?              �?      @              :@     r@      $@     �J@      @      E@              3@      @      7@      @      *@       @      �?              �?       @              �?      (@              "@      �?      @              @      �?                      $@      @      &@      @              �?      &@      �?       @               @      �?                      "@      0@     �m@      @      c@             �H@      @      Z@      @     �F@      @      >@              *@      @      1@       @              @      1@       @      (@       @      "@       @      @              @       @                      @              @      @      @       @      @       @       @               @       @                      @      �?                      .@             �M@      "@     �T@       @      @      �?              �?      @              @      �?              @     �S@      @      I@      �?              @      I@              0@      @      A@      @      @      @      �?      @                      �?              @      @      =@      �?      =@              :@      �?      @      �?                      @       @                      =@     �q@      T@     �M@      L@      L@      F@     �I@      9@      @      *@      �?      *@      �?      �?              �?      �?                      (@       @              H@      (@      2@      �?      @      �?       @      �?      �?      �?      �?                      �?      �?              �?              .@              >@      &@      2@      �?       @      �?       @                      �?      0@              (@      $@      (@      @      �?      @      �?                      @      &@       @      &@                       @              @      @      3@       @      2@       @      &@      �?      "@              "@      �?              �?       @               @      �?                      @      @      �?              �?      @              @      (@      �?      (@      �?      @      �?                      @              @       @             �l@      8@     �l@      3@      @       @              @      @      @      @      �?      @                      �?              @     �k@      &@      :@      @              @      :@      @      8@               @      @       @                      @     �h@      @     `h@      @     @h@       @     `d@              ?@       @               @      ?@              �?      �?      �?                      �?       @       @       @                       @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��-hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�BX7         z                    �?�6𿸴�?:           ��@                           _@�e�,��?K           ��@                           �?6YE�t�?0            �P@                          P`@���|���?             6@                           �I@d}h���?             ,@                           `@      �?             @������������������������       �                      @������������������������       �                      @	       
                    �?ףp=
�?             $@������������������������       �                     @                          �`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @              
             �?      �?              @������������������������       �                     @������������������������       �                     @                           �?���7�?              F@������������������������       �                     B@                          @c@      �?              @������������������������       �                     @              	          `ff@�q�q�?             @������������������������       �                     �?������������������������       �                      @       G       
             �?
��^���?           }@                            �?��R���?h            �e@                          �b@r�q��?             H@                           �?Du9iH��?            �E@              	          `ff@��Y��]�?            �D@������������������������       �                     D@������������������������       �                     �?������������������������       �                      @������������������������       �                     @!       ,                    �?x�����?M             _@"       #                    �?Hث3���?            �C@������������������������       �        
             ,@$       %                    �L@�+e�X�?             9@������������������������       �                     *@&       '                   �a@      �?             (@������������������������       �                     @(       +                    �N@      �?              @)       *       	          ���@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @-       .       	          833�?������?4            @U@������������������������       �                     @@/       @                   d@䯦s#�?!            �J@0       ;                    �N@>A�F<�?             C@1       2       	          833�?<���D�?            �@@������������������������       �                      @3       :                    �?`Jj��?             ?@4       5                   �Q@�t����?             1@������������������������       �                     �?6       7                   hq@      �?
             0@������������������������       �                     *@8       9                   @]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             ,@<       =                   @_@���Q��?             @������������������������       �                     �?>       ?                    �P@      �?             @������������������������       �                     @������������������������       �                     �?A       B                    @G@�r����?             .@������������������������       �                     @C       F                   0m@      �?              @D       E                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @H       c                    @L@��P��?�            Pr@I       b                   h@�?�|�?�            �k@J       M                   @c@�:�h���?�            �k@K       L                    �?      �?              @������������������������       �                     �?������������������������       �                     �?N       [                   @\@�HGݐ\�?�            `k@O       R                   �e@l��\��?             A@P       Q                    @F@�q�q�?             @������������������������       �                     �?������������������������       �                      @S       Z       	          ����?`Jj��?             ?@T       U                    �E@�8��8��?             8@������������������������       �                     &@V       Y                   Pc@8�Z$���?             *@W       X                   �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     "@������������������������       �                     @\       a                    �? S5W�?n             g@]       ^       	            �?P�Lt�<�?             C@������������������������       �                     ?@_       `       	          ����?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �        W            `b@������������������������       �                     �?d       u                    �N@\�CX�?)            �Q@e       f                    i@X�Cc�?             E@������������������������       �                     &@g       l                   �a@�g�y��?             ?@h       k                    �?�8��8��?             (@i       j                    @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @m       t                    �?�d�����?             3@n       s                   0f@      �?
             0@o       r                    �?��S�ۿ?	             .@p       q       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?������������������������       �                     @v       w                   p@XB���?             =@������������������������       �        
             .@x       y                    �?@4և���?	             ,@������������������������       �                     �?������������������������       �                     *@{       �       
             �?Pp	~86�?�            0x@|       �                    �?�������?�            `t@}       �                   �Z@H�̱���?�            @o@~       �                   �Y@և���X�?             @       �                   0a@z�G�z�?             @������������������������       �                     @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �b@�g�H��?�            `n@�       �                    �?�Ȍ���?�            �l@�       �                    �?؇���X�?             5@�       �                   h@�KM�]�?             3@������������������������       �                     �?�       �       	          ����?�X�<ݺ?             2@�       �                    @J@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@�       �                    `@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �R@��+��?�            �i@�       �                    �?�:���ΰ?            �i@�       �                    �D@@�E�x�?Z            `b@�       �                    `@ףp=
�?             $@�       �       	          ����?�q�q�?             @������������������������       �                     �?�       �                    e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �_@ ���v�?S             a@�       �       	          hff�?����D��?<            @W@�       �                    �?$�q-�?
             *@�       �                    @O@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @�       �                   0i@@�z�G�?2             T@�       �                    \@Pa�	�?            �@@�       �       
             �?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@������������������������       �                    �G@������������������������       �                     F@�       �                   `\@ ,��-�?%            �M@�       �       
             �?d}h���?             ,@������������������������       �                     �?�       �                    �L@�θ�?
             *@�       �                    Z@���Q��?             @�       �                    @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       
             �?����?�?            �F@������������������������       �                     &@�       �                   �]@г�wY;�?             A@�       �                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @@������������������������       �                     �?�       �                    �?�r����?	             .@�       �                   pk@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	          `ff�?�8��8��?             (@������������������������       �                     "@�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �s@���y4F�?*             S@�       �                   �[@�ˡ�5��?(            �Q@�       �                    �H@����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �J@     ��?"             P@�       �                    �I@�q�q�?             .@�       �       	          033�?�θ�?             *@������������������������       �                     @�       �                   �l@      �?             @�       �                    �G@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �       	          ����?@9G��?            �H@�       �                   @e@@4և���?             <@�       �                    �? 7���B�?             ;@�       �                    n@      �?	             0@������������������������       �                     &@�       �                   o@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                     �?������������������������       �        
             5@�       �                   �^@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��7��?)            �N@�       �                    @N@�T|n�q�?            �E@�       �       	             �?��a�n`�?             ?@�       �                   �a@X�<ݚ�?             "@�       �                   �`@�q�q�?             @������������������������       �                      @�       �                   `k@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	          `ff�?�C��2(�?             6@�       �                    @M@P���Q�?             4@������������������������       �                     *@�       �                    �?؇���X�?             @�       �       	          033�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�       �                   pa@�����H�?             2@������������������������       �                      @�       �                   @b@z�G�z�?             $@������������������������       �                      @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     p@     �v@     `e@      $@      L@       @      ,@      @      &@       @       @       @                       @      �?      "@              @      �?      @      �?                      @      @      @              @      @               @      E@              B@       @      @              @       @      �?              �?       @             �u@     �\@     �S@     @W@      D@       @      D@      @      D@      �?      D@                      �?               @              @     �C@     @U@      3@      4@              ,@      3@      @      *@              @      @              @      @       @      �?       @               @      �?              @              4@     @P@              @@      4@     �@@      @      ?@      @      =@       @               @      =@       @      .@      �?              �?      .@              *@      �?       @               @      �?                      ,@      @       @              �?      @      �?      @                      �?      *@       @      @              @       @      �?       @               @      �?              @             �p@      6@      k@      @      k@      @      �?      �?              �?      �?             �j@      @      ?@      @       @      �?              �?       @              =@       @      6@       @      &@              &@       @       @       @       @                       @      "@              @              g@      �?     �B@      �?      ?@              @      �?              �?      @             `b@                      �?     �K@      0@      ;@      .@      &@              0@      .@      &@      �?      @      �?      @                      �?      @              @      ,@       @      ,@      �?      ,@      �?      �?              �?      �?                      *@      �?              @              <@      �?      .@              *@      �?              �?      *@             �K@     �t@      @@     `r@      0@     @m@      @      @      �?      @              @      �?      �?              �?      �?               @              *@     �l@      &@      k@      @      2@       @      1@      �?              �?      1@      �?      @      �?                      @              ,@      �?      �?              �?      �?               @     �h@      @     �h@      @      b@      �?      "@      �?       @              �?      �?      �?              �?      �?                      @       @     �`@       @     �V@      �?      (@      �?      "@              "@      �?                      @      �?     �S@      �?      @@      �?      @              @      �?                      ;@             �G@              F@      @     �K@      @      &@              �?      @      $@      @       @      �?       @               @      �?               @                       @      �?      F@              &@      �?     �@@      �?      �?      �?                      �?              @@      �?               @      *@      �?       @               @      �?              �?      &@              "@      �?       @      �?                       @      0@      N@      (@     �M@      @       @               @      @              @     �L@      @      $@      @      $@              @      @      @      @      �?      @                      �?               @       @               @     �G@       @      :@      �?      :@      �?      .@              &@      �?      @      �?                      @              &@      �?                      5@      @      �?      @                      �?      7@      C@      @      B@      @      8@      @      @       @      @               @       @       @               @       @              @               @      4@      �?      3@              *@      �?      @      �?       @               @      �?                      @      �?      �?              �?      �?                      (@      0@       @       @               @       @               @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�m7hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKㅔh~�B�1         �                    �?@���u�?>           ��@       !                    �?�$xV{�?9           0�@              	          033�?:�1�(��?2            @U@                          �b@ �o_��?             I@                           a@\X��t�?             7@                          a@؇���X�?	             ,@������������������������       �                     $@              
             �?      �?             @	       
                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?                          �`@�����H�?             "@                          @e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                           \@PN��T'�?             ;@������������������������       �                     �?                           @P@ȵHPS!�?             :@                           �? �q�q�?             8@              
             �?�C��2(�?             &@������������������������       �                     @                          �d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@������������������������       �                      @                            ]@ >�֕�?            �A@                           k@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @@"       Y       
             �?��!�?           {@#       V                    �?T�	�S�?�             u@$       U                   �e@�θV�?�            �i@%       *                    �?l��\��?�            �i@&       '                    `P@      �?             @@������������������������       �                     >@(       )                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?+       T                   �a@��0��?m            �e@,       M                   (q@�0&���?S            @_@-       J                    c@�!��U��??            �W@.       I       	          ����?�k��?:            @V@/       4                    @K@�z�6�?)             O@0       1                   Pm@���7�?             6@������������������������       �                     2@2       3                    `@      �?             @������������������������       �                     @������������������������       �                     �?5       6       	          ����?�z�G��?             D@������������������������       �                     &@7       :       	             �?�f7�z�?             =@8       9                    X@r�q��?             @������������������������       �                     �?������������������������       �                     @;       D                    �L@8����?             7@<       C                   �`@���Q��?             $@=       >       	          ����?      �?              @������������������������       �                     @?       @                    @L@���Q��?             @������������������������       �                     �?A       B                    ^@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @E       H       
             �?$�q-�?             *@F       G                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     ;@K       L                    @L@      �?             @������������������������       �                     @������������������������       �                     @N       S                    �?(;L]n�?             >@O       P                    �G@      �?              @������������������������       �                     @Q       R       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@������������������������       �                    �G@������������������������       �                     @W       X                    �R@ g�yB�?E             `@������������������������       �        D            �_@������������������������       �                      @Z       q       	          833�?�E���?@            @X@[       f                   �a@��C���?"            �G@\       ]       	             �PN��T'�?             ;@������������������������       �                     �?^       e                   �`@ȵHPS!�?             :@_       `                    W@d}h���?             ,@������������������������       �                      @a       d                    �?�8��8��?	             (@b       c       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     (@g       p                   Xs@      �?             4@h       i                   �d@r�q��?             2@������������������������       �                      @j       k                    @C@�z�G��?             $@������������������������       �                      @l       m                     K@      �?              @������������������������       �                     @n       o                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @r              	          033�?�J�4�?             I@s       ~                    �?������?            �D@t       }                   �s@���y4F�?             3@u       x                    @F@�t����?             1@v       w                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?y       |       	          ����?@4և���?	             ,@z       {                    ]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                      @������������������������       �                     6@�       �                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�       �       
             �?���Q8�?            y@�       �       	          ����?��Y���?c            �c@�       �       
             �?��2(&�?             F@������������������������       �                      @�       �                   @`@�����?             E@������������������������       �                     :@�       �                   �`@      �?
             0@������������������������       �                      @�       �                   �j@؇���X�?	             ,@�       �                   �f@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �N@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?�s��:��?I            �\@�       �                   `\@��j��?1            @S@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                   d@�û��|�?,            @Q@�       �                     J@��B����?"             J@�       �                    �?�C��2(�?             &@�       �       	              @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    `@��]�T��?            �D@�       �       	          033�?��
ц��?	             *@�       �                   @[@�q�q�?             "@������������������������       �                     �?�       �       	             �?      �?              @�       �                    �?      �?             @�       �                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?����X�?             <@�       �       
             �?r�q��?             (@������������������������       �                     @�       �                   �n@����X�?             @�       �                   �c@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    @      �?             0@�       �                    �K@      �?             (@������������������������       �                      @�       �                   �^@�z�G��?             $@�       �                     R@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    a@�t����?
             1@������������������������       �        	             .@������������������������       �                      @�       �                   �^@���@��?            �B@�       �       
             �?X�<ݚ�?             "@������������������������       �                     @�       �                   `c@r�q��?             @�       �                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �`@ �Cc}�?             <@������������������������       �                     5@�       �                   �o@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                   �g@��a��?�            @n@�       �       	          ���@x�e�� �?�             n@�       �       	            �?(�5�f��?�            �m@�       �                   @[@���ۮ��?�            �h@�       �                   0n@�����H�?
             2@������������������������       �                     .@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        z            `f@�       �                    @z�G�z�?             D@�       �                   �e@��hJ,�?             A@������������������������       �                     @�       �       	          ����?`Jj��?             ?@�       �                   �p@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     8@�       �                    a@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�B0       �w@     ��@     @X@     Pz@      C@     �G@      B@      ,@      *@      $@      (@       @      $@               @       @      �?       @               @      �?              �?              �?       @      �?      @              @      �?                      @      7@      @              �?      7@      @      7@      �?      $@      �?      @              @      �?      @                      �?      *@                       @       @     �@@       @      �?       @                      �?              @@     �M@     `w@      7@     �s@      5@     @g@      2@     @g@      �?      ?@              >@      �?      �?              �?      �?              1@     `c@      1@      [@      0@     �S@      *@      S@      *@     �H@      �?      5@              2@      �?      @              @      �?              (@      <@              &@      (@      1@      @      �?              �?      @              @      0@      @      @      @       @      @              @       @              �?      @      �?      @                      �?               @      �?      (@      �?       @      �?                       @              $@              ;@      @      @              @      @              �?      =@      �?      @              @      �?      �?              �?      �?                      6@             �G@      @               @     �_@             �_@       @              B@     �N@      <@      3@      7@      @              �?      7@      @      &@      @               @      &@      �?      �?      �?      �?                      �?      $@              (@              @      .@      @      .@               @      @      @       @              �?      @              @      �?      �?              �?      �?               @               @      E@      @     �B@      @      .@       @      .@      �?       @               @      �?              �?      *@      �?      �?              �?      �?                      (@       @                      6@      @      @      @                      @     �q@     �\@     �L@     @Y@      @      C@       @              @      C@              :@      @      (@       @               @      (@      �?       @               @      �?              �?      $@              $@      �?             �I@     �O@     �E@      A@      �?      @      �?                      @      E@      ;@      ;@      9@      �?      $@      �?       @      �?                       @               @      :@      .@      @      @      @      @              �?      @       @       @       @       @      �?       @                      �?              �?      @                      @      4@       @      $@       @      @              @       @      @      �?              �?      @                      �?      $@      @      "@      @       @              @      @       @      @              @       @              @              �?      @      �?                      @      .@       @      .@                       @       @      =@      @      @              @      @      �?       @      �?       @                      �?      @              @      9@              5@      @      @      @                      @     �l@      ,@     �l@      *@     �l@      "@     `h@       @      0@       @      .@              �?       @      �?                       @     `f@             �@@      @      =@      @              @      =@       @      @       @               @      @              8@              @       @               @      @                      @              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�2�hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKh~�BH4         �       
             �?���ƒ�?>           ��@       I                    �?��yF��?G           p�@       @                    �?L
e��?�            �i@              	          ����?b��H���?Z            �b@                           �?�2����?             �K@������������������������       �                     :@                           a@8^s]e�?             =@       	                    �?�8��8��?             (@������������������������       �                      @
                           �K@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?                           �?��.k���?             1@                           �J@�q�q�?             "@������������������������       �                     @                          p@���Q��?             @������������������������       �                     @������������������������       �                      @                           g@      �?              @              
             �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?       7       	          033�?ܐ҆��?:            @W@       "                   �b@�c�Α�?$             M@                          �n@ףp=
�?             >@������������������������       �        	             0@                           �?d}h���?             ,@������������������������       �                     "@                          `@���Q��?             @������������������������       �                      @        !                   �q@�q�q�?             @������������������������       �                     �?������������������������       �                      @#       $                   �b@���>4��?             <@������������������������       �                     @%       &                   �K@���Q��?             9@������������������������       �                      @'       (       
             �?�LQ�1	�?             7@������������������������       �                     @)       0                   �^@      �?             4@*       /                    �?$�q-�?             *@+       ,                    @I@�q�q�?             @������������������������       �                     �?-       .                     O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@1       2                    �I@և���X�?             @������������������������       �                     @3       4       	          ����?      �?             @������������������������       �                      @5       6                    �?      �?              @������������������������       �                     �?������������������������       �                     �?8       =                    �?(N:!���?            �A@9       <                   �u@���!pc�?             &@:       ;                    �O@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @>       ?                   �d@ �q�q�?             8@������������������������       �                     7@������������������������       �                     �?A       H                   �g@�j��b�?&            �M@B       C                    �?l�b�G��?%            �L@������������������������       �                     D@D       E                   �a@������?             1@������������������������       �                      @F       G                    d@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @J       O                   �Z@0`%w�?�            �s@K       N                    �?և���X�?             @L       M                   Pa@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @P       W                   Pe@��T����?�            �s@Q       V                    I@`���i��?6             V@R       S                   0a@�?�|�?-            �R@������������������������       �        (            �P@T       U                    �?����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             ,@X       �                   �b@���>4��?�             l@Y       �                    @T�y���?�            `j@Z                          ``@�R��ݽ?�             j@[       `                    �?H��?"�?2             U@\       ]                    @P@���N8�?             5@������������������������       �        
             2@^       _                    �P@�q�q�?             @������������������������       �                     �?������������������������       �                      @a       d                   �f@��d��?%            �O@b       c                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @e       t                   `\@�r����?#             N@f       s       	             @�q�q�?             2@g       p                   �Z@      �?
             0@h       m                    �?8�Z$���?             *@i       j                    _@ףp=
�?             $@������������������������       �                     @k       l       	          433�?      �?             @������������������������       �                     �?������������������������       �                     @n       o                    @K@�q�q�?             @������������������������       �                      @������������������������       �                     �?q       r                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @u       ~                    ^@���N8�?             E@v       }                    �?8�Z$���?             *@w       x                    @M@�8��8��?             (@������������������������       �                     @y       z       	             �?z�G�z�?             @������������������������       �                     �?{       |                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     =@�       �                    �?@�n�1�?P            @_@�       �                   �b@�D�e���?7            @U@������������������������       �                     G@�       �                    @F@�7��?            �C@������������������������       �                     �?�       �                    �?P�Lt�<�?             C@������������������������       �                     8@�       �                    �Q@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                     D@������������������������       �                      @�       �                    �?�n_Y�K�?	             *@�       �                    @O@���!pc�?             &@�       �                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    �?�ME6���?�            �x@�       �                   @E@dq5n��?�            �u@�       �                    �?��.k���?             A@������������������������       �                     �?�       �                   �[@�'�=z��?            �@@�       �                   �_@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?X�<ݚ�?             ;@�       �                   �\@r�q��?
             (@������������������������       �                      @������������������������       �        	             $@�       �                    �?�r����?	             .@�       �                    `Q@@4և���?             ,@������������������������       �                     &@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    �L@l,��?�            `s@�       �                   �k@8������?�            �o@�       �                    �?P�c0"�?A            @Z@�       �       	             �?��:�-�?=            @Y@������������������������       �        7            �V@�       �                    �?z�G�z�?             $@�       �                    _@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @�       �                   �i@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �f@��'#��?X            �b@�       �                   @[@�w�uz
�?U            �a@�       �                    �?      �?              @������������������������       �                     @������������������������       �                     @�       �                    �?����?�?R            �`@�       �                    �?؇���X�?             5@������������������������       �                     (@�       �                   @_@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �        F            �\@�       �                    �C@���Q��?             @������������������������       �                     �?�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �b@�k�'7��?&            �L@�       �       	          033@ >�֕�?            �A@�       �                    ]@г�wY;�?             A@�       �                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @@������������������������       �                     �?�       �                   �`@���|���?             6@�       �                    �M@r�q��?             @������������������������       �                     @�       �                   �c@�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    b@     ��?	             0@�       �                   pr@�z�G��?             $@������������������������       �                     @�       �                   �c@      �?             @�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?�q�q�?!             H@�       �       	          ����?R���Q�?             D@�       �                    �?ҳ�wY;�?             1@�       �                    n@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�q�q�?             (@�       �                   �`@�z�G��?             $@�       �                    @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     7@������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       `y@      �@     @V@     P{@     �N@     @b@     �K@     @W@      "@      G@              :@      "@      4@      �?      &@               @      �?      "@              "@      �?               @      "@      @      @      @               @      @              @       @               @      @      �?      @      �?                      @      �?              G@     �G@      E@      0@      ;@      @      0@              &@      @      "@               @      @               @       @      �?              �?       @              .@      *@              @      .@      $@               @      .@       @              @      .@      @      (@      �?       @      �?      �?              �?      �?              �?      �?              $@              @      @              @      @      �?       @              �?      �?      �?                      �?      @      ?@      @       @      @      @              @      @                      @      �?      7@              7@      �?              @     �J@      @     �J@              D@      @      *@               @      @      @      @                      @       @              <@     0r@      @      @      @       @               @      @                       @      9@     �q@       @     �U@       @      R@             �P@       @      @              @       @                      ,@      7@      i@      .@     �h@      *@     �h@      &@     @R@      �?      4@              2@      �?       @      �?                       @      $@     �J@       @      �?              �?       @               @      J@      @      (@      @      (@       @      &@      �?      "@              @      �?      @      �?                      @      �?       @               @      �?               @      �?       @                      �?       @               @      D@       @      &@      �?      &@              @      �?      @              �?      �?      @      �?                      @      �?                      =@       @     �^@       @     �T@              G@       @     �B@      �?              �?     �B@              8@      �?      *@              *@      �?                      D@       @               @      @       @      @       @       @       @                       @              �?               @     �s@     �R@     �r@     �D@      0@      2@              �?      0@      1@      �?      @              @      �?              .@      (@       @      $@       @                      $@      *@       @      *@      �?      &@               @      �?       @                      �?              �?     �q@      7@      n@      *@     �Y@       @     �X@       @     �V@               @       @      �?      �?              �?      �?              @      �?      @              @      �?      @                      �?      @              a@      &@     �`@       @      @      @      @                      @     �`@      @      2@      @      (@              @      @              @      @             �\@               @      @      �?              �?      @      �?                      @     �G@      $@     �@@       @     �@@      �?      �?      �?              �?      �?              @@                      �?      ,@       @      �?      @              @      �?       @              �?      �?      �?              �?      �?              *@      @      @      @      @              �?      @      �?      �?              �?      �?                       @      @              ,@      A@      @      A@      @      &@      �?      @      �?                      @      @      @      @      @       @      �?              �?       @              �?      @      �?                      @       @                      7@       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��^ZhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �                    �?��+�?T           ��@       O                    �J@��M�
��?D           p@       ,       
             �?n,
#9�?�            �j@                           �?$s��O�?[            �a@                          �e@Hm_!'1�?            �H@              	          ����?`�q�0ܴ?            �G@������������������������       �                     A@       	                   hp@8�Z$���?             *@������������������������       �                     $@
                          �u@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                           �?؇���X�?=            �V@                          �`@��S���?             .@              	          ����?�<ݚ�?             "@                          �[@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @       %                   pa@`-�I�w�?6             S@               	             @���U�?)            �L@                           �D@ pƵHP�?%             J@                           e@�C��2(�?	             &@������������������������       �                     @              
             �?z�G�z�?             @������������������������       �                     �?                           `@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �D@!       "                   �Z@z�G�z�?             @������������������������       �                     @#       $                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?&       +                    @J@�S����?             3@'       *                   �b@�����H�?             2@(       )                   �\@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     &@������������������������       �                     �?-       <                   �a@l�;�	�?4            �R@.       1                    �?\-��p�?             =@/       0                   �a@���Q��?             @������������������������       �                     @������������������������       �                      @2       3                   �\@�8��8��?             8@������������������������       �                     @4       5                   �^@�t����?             1@������������������������       �                     @6       9                    �?"pc�
�?
             &@7       8                    P@�����H�?             "@������������������������       �                     �?������������������������       �                      @:       ;       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?=       >                    �?��c:�?             G@������������������������       �                      @?       N                   �f@p9W��S�?             C@@       M                    �?H�V�e��?             A@A       H                   �`@R�}e�.�?             :@B       C                   d@      �?             0@������������������������       �                     &@D       E                    �?z�G�z�?             @������������������������       �                     �?F       G       	             �?      �?             @������������������������       �                     �?������������������������       �                     @I       J                    �D@���Q��?             $@������������������������       �                      @K       L                    �?      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @P       u       
             �?���Hx�?�             r@Q       t                   {@�NI���?�             m@R       q                   �c@��F�M�?�            �l@S       Z                    �?�'B���?�            �k@T       Y                    `@z�G�z�?             9@U       V                   �`@�eP*L��?	             &@������������������������       �                     @W       X                    _@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             ,@[       \                    �?��~F�<�?z            �h@������������������������       �                     A@]       p                   �_@��w#'�?f            `d@^       o                    �R@ЮN
��?G            @\@_       l                   `_@�v�ɱ?F            �[@`       k       	          ����?P�c0"�?C            @Z@a       j                    `@      �?-             P@b       g       	          033�? 	��p�?             =@c       d       	          ����? ��WV�?             :@������������������������       �        	             ,@e       f                   �_@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?h       i                    �M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                    �A@������������������������       �                    �D@m       n                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     I@r       s                   @d@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @v       y                    �L@4և����?"             L@w       x                    �?      �?              @������������������������       �                     @������������������������       �                     @z       �                   Pl@r�q��?             H@{       �                   �a@�X����?             6@|       �       	          033�?      �?             0@}       ~                    �?��S�ۿ?
             .@������������������������       �                     (@       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �e@ ��WV�?             :@������������������������       �                     9@������������������������       �                     �?�       �       
             �?�Kc��-�?           �y@�       �                    �?d��J_��?f            `c@�       �       
             �?z�J��?B            �W@�       �                   �]@�r����?
             .@������������������������       �                      @������������������������       �                     *@�       �                    �?���;+"�?8            �S@�       �       	          ���ٿ��>4և�?             <@������������������������       �                     @�       �                    @L@`�Q��?             9@������������������������       �                     "@�       �                   0b@      �?             0@�       �                    �?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�       �                    �?؇���X�?             @�       �                   pk@r�q��?             @�       �                    `Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    �?�\�u��?%            �I@�       �                    �?�G�z��?             4@�       �                   �b@     ��?             0@�       �       	          ����?d}h���?
             ,@�       �                    �?�q�q�?             "@�       �       	             �?      �?             @������������������������       �                     �?�       �                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   0n@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   0a@�חF�P�?             ?@�       �                   �`@�E��ӭ�?             2@�       �                    �?z�G�z�?             .@�       �                    �K@�C��2(�?	             &@������������������������       �                     "@�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   `b@      �?             @������������������������       �                     �?�       �       	          `ff@�q�q�?             @������������������������       �                     �?�       �       	          `ff@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             *@�       �                   Pe@`��:�?$            �N@������������������������       �                     .@�       �                    c@��+7��?             G@�       �                    �J@z�G�z�?             D@������������������������       �                     �?�       �                   �\@8�Z$���?            �C@������������������������       �                     @�       �                   �`@г�wY;�?             A@�       �                   �[@�����H�?             "@������������������������       �                     @�       �                   �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     9@�       �       	          ���@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?��a�!��?�            @p@�       �                    @G@`�q��־?�             m@������������������������       �        @            @Y@�       �                    f@�Ra����?W            �`@�       �                    �?ףp=
�?V            @`@�       �       	          033@POͳF��?P            �]@�       �                     R@ج��w�?O            �\@�       �                   �l@l�b�G��?N            �\@�       �                    �H@��<b�ƥ?              G@�       �                   P`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �E@�       �       	          pff�?ДX��?.             Q@�       �                     L@���V��?            �F@�       �                    �?�>����?             ;@������������������������       �                     3@�       �                   �c@      �?              @�       �                    �?      �?             @������������������������       �                     �?�       �                   �n@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �m@�E��ӭ�?             2@������������������������       �                      @�       �                   �c@     ��?             0@�       �                    �L@�r����?
             .@������������������������       �                     �?�       �                   �c@@4և���?	             ,@�       �                   pa@؇���X�?             @������������������������       �                      @�       �       	          ����?z�G�z�?             @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     7@������������������������       �                     �?������������������������       �                     @������������������������       �                     &@������������������������       �                      @�             	          033�?������?             ;@                         Hs@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?                         �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�t�b�*     h�h(h+K ��h-��R�(KMKK��h_�BP       x@     ��@     @V@     �y@     �N@     @c@      1@     �^@      @     �F@       @     �F@              A@       @      &@              $@       @      �?       @                      �?       @              *@     �S@       @      @       @      @       @       @               @       @                      @      @              @     �Q@       @     �K@      �?     �I@      �?      $@              @      �?      @              �?      �?      @      �?                      @             �D@      �?      @              @      �?      �?              �?      �?              @      0@       @      0@       @      @       @                      @              &@      �?              F@      ?@      9@      @      @       @      @                       @      6@       @      @              .@       @      @              "@       @       @      �?              �?       @              �?      �?      �?                      �?      3@      ;@       @              &@      ;@      @      ;@      @      3@      �?      .@              &@      �?      @              �?      �?      @      �?                      @      @      @               @      @       @      @                       @               @      @              <@     @p@      .@      k@      *@      k@      &@     `j@      @      4@      @      @      @              �?      @              @      �?                      ,@      @     �g@              A@      @     �c@      @     �Z@      @     �Z@       @     �Y@       @      O@       @      ;@      �?      9@              ,@      �?      &@              &@      �?              �?       @               @      �?                     �A@             �D@       @      @       @                      @       @                      I@       @      @       @                      @       @              *@     �E@      @      @      @                      @       @      D@      @      .@       @      ,@      �?      ,@              (@      �?       @      �?                       @      �?              @      �?      @                      �?      �?      9@              9@      �?             �r@     �]@      M@     @X@      G@      H@      *@       @               @      *@             �@@      G@      1@      &@              @      1@       @      "@               @       @       @      @       @                      @      @      �?      @      �?       @      �?              �?       @              @              �?              0@     �A@      &@      "@      &@      @      &@      @      @      @       @       @      �?              �?       @               @      �?              @      �?      @                      �?      @                       @              @      @      :@      @      *@      @      (@      �?      $@              "@      �?      �?      �?                      �?       @       @              �?       @      �?      �?              �?      �?              �?      �?               @      �?       @                      �?              *@      (@     �H@              .@      (@      A@      @     �@@      �?              @     �@@      @              �?     �@@      �?       @              @      �?      @              @      �?                      9@      @      �?      @                      �?     �m@      6@     @k@      .@     @Y@             @]@      .@     @]@      *@     �Z@      *@     �Z@      "@     �Z@       @     �F@      �?       @      �?              �?       @             �E@             �N@      @      C@      @      9@       @      3@              @       @       @       @      �?              �?       @               @      �?              @              *@      @               @      *@      @      *@       @              �?      *@      �?      @      �?       @              @      �?      �?      �?      �?                      �?      @              @                      �?      7@                      �?              @      &@                       @      4@      @      3@      �?      3@                      �?      �?      @      �?                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJтhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKׅ�h~�B/         �                    �?���3L�?7           ��@       1                    �?��+��?�           ��@                           �?z�G�z�?i            @e@              
             �?�θV�?S            @a@                           �?P����?             C@                           @E@D�n�3�?             3@������������������������       �                      @       	                   @d@��.k���?             1@������������������������       �                      @
                           b@���Q��?             .@              	          ����?�q�q�?             "@                          Pb@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @              	          ����?�KM�]�?             3@                          `X@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     &@                           T@ �ׁsF�?9             Y@������������������������       �                     �?������������������������       �        8            �X@       ,                    �?      �?             @@       %                   �`@�GN�z�?             6@                            b@      �?              @              	          433�?z�G�z�?             @������������������������       �                      @              	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @!       "                   �d@�q�q�?             @������������������������       �                     �?#       $                     L@      �?              @������������������������       �                     �?������������������������       �                     �?&       '                    @H@؇���X�?	             ,@������������������������       �                     �?(       )       	          ����?$�q-�?             *@������������������������       �                     &@*       +                   Pc@      �?              @������������������������       �                     �?������������������������       �                     �?-       .                   @_@�z�G��?             $@������������������������       �                     @/       0       	             �?      �?             @������������������������       �                     @������������������������       �                     @2       m       	          pff�?(�q;Y9�?G           ��@3       <                   @E@8����;�?�            �r@4       5       
             �?������?            �D@������������������������       �                     >@6       ;       	            �?���|���?             &@7       8                   �Y@և���X�?             @������������������������       �                      @9       :                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @=       L       
             �?P�>�,��?�            p@>       A       	          ����?�㙢�c�?&            @Q@?       @                    g@ �Jj�G�?            �K@������������������������       �                     K@������������������������       �                     �?B       G                    �?d}h���?             ,@C       F                   �i@ףp=
�?             $@D       E                    @N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @H       I                   �^@      �?             @������������������������       �                     �?J       K                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @M       Z                    �I@�*/�8V�?t            �g@N       S                    �?Xc!J�ƴ?H            �]@O       R                    e@z�G�z�?             .@P       Q                   �`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@T       Y                   @[@p� V�?=            �Y@U       V                    �E@"pc�
�?             &@������������������������       �                     @W       X                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        8             W@[       h                   pc@d}h���?,            �Q@\       e                    @Hm_!'1�?             �H@]       b                   �o@=QcG��?            �G@^       _                    �?P�Lt�<�?             C@������������������������       �                    �A@`       a       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?c       d                   Xp@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @f       g                   ``@      �?              @������������������������       �                     �?������������������������       �                     �?i       j                    �?�G��l��?             5@������������������������       �                      @k       l                   �f@�θ�?             *@������������������������       �                     $@������������������������       �                     @n       �       	          033�?�Y	��o�?�            `m@o       x                    _@��xKm�?P            �_@p       q                    �?h㱪��?!            �K@������������������������       �                    �B@r       s                   �f@�����H�?             2@������������������������       �                      @t       w                    �?z�G�z�?             $@u       v                   Pk@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @y       �                   �b@F��ӭ��?/             R@z       {       	          `ff�?F�����?            �F@������������������������       �                     @|       �                    b@H�z�G�?             D@}       �                    �?�q�q�?            �@@~       �                   �_@R���Q�?             4@       �                   �^@���Q��?             @�       �                   l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   �[@��S�ۿ?             .@�       �                   �j@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             (@�       �                   �`@�n_Y�K�?             *@�       �                   @m@���!pc�?             &@������������������������       �                     @�       �                    �K@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �_@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    @�q�q�?             ;@�       �                    �?��+7��?             7@�       �                   m@      �?
             0@�       �                   �i@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     (@�       �                    �?և���X�?             @������������������������       �                     @������������������������       �                     @�       �       
             �?      �?             @������������������������       �                     �?������������������������       �                     @�       �       
             �? 7���B�?C             [@�       �       	          `ff@��:�-�?>            @Y@�       �                   �Z@�eGk�T�?9            �W@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        7             W@�       �                   �a@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?����X�?             @�       �                    �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?(L���?�            �j@�       �                    �? �й���?_            @b@�       �                    @J@��ɉ�?)            @P@�       �       	          ����?�����H�?             2@������������������������       �        	             &@�       �       
             �?����X�?             @������������������������       �                     @�       �                   �b@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                    �G@������������������������       �        6            @T@�       �                    �?��x�5��?(            @Q@�       �       
             �?�>$�*��?            �D@�       �                   ``@�q�q�?             2@�       �                   @c@      �?              @������������������������       �                     @������������������������       �                     @�       �                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                   �U@��+7��?             7@������������������������       �                     @�       �                   xs@R���Q�?             4@�       �                   �`@�X�<ݺ?             2@�       �                    �O@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             ,@������������������������       �                      @�       �                   �Z@�>4և��?             <@������������������������       �                     @�       �                    �N@HP�s��?             9@�       �                    �?8�Z$���?             *@�       �                     M@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   0b@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     (@�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp       px@     x�@     �v@     `u@      a@      A@      _@      ,@      9@      *@       @      &@               @       @      "@       @              @      "@      @      @       @      @       @                      @      @                      @      1@       @      @       @               @      @              &@             �X@      �?              �?     �X@              (@      4@      @      1@      @      @      �?      @               @      �?       @      �?                       @       @      �?      �?              �?      �?              �?      �?               @      (@      �?              �?      (@              &@      �?      �?      �?                      �?      @      @      @              @      @              @      @              l@     @s@      g@     �\@      @     �B@              >@      @      @      @      @               @      @      �?      @                      �?              @     �f@     @S@      (@     �L@      �?      K@              K@      �?              &@      @      "@      �?      �?      �?      �?                      �?       @               @       @      �?              �?       @      �?                       @      e@      4@     @\@      @      (@      @      �?      @              @      �?              &@             @Y@       @      "@       @      @              @       @      @                       @      W@             �K@      .@     �F@      @      F@      @     �B@      �?     �A@               @      �?       @                      �?      @       @               @      @              �?      �?              �?      �?              $@      &@               @      $@      @      $@                      @     �D@     @h@     �B@     �V@       @     �J@             �B@       @      0@               @       @       @       @      @       @                      @               @     �A@     �B@      1@      <@              @      1@      7@      &@      6@      @      1@       @      @       @      �?       @                      �?               @      �?      ,@      �?       @               @      �?                      (@       @      @       @      @      @              �?      @              @      �?                       @      @      �?              �?      @              2@      "@      1@      @      ,@       @       @       @       @                       @      (@              @      @              @      @              �?      @      �?                      @      @      Z@       @     �X@      �?     �W@      �?       @      �?                       @              W@      �?      @              @      �?               @      @       @      �?              �?       @                      @      >@      g@       @      b@       @     �O@       @      0@              &@       @      @              @       @       @       @                       @             �G@             @T@      <@     �D@      7@      2@      @      (@      @      @              @      @              �?      "@      �?                      "@      1@      @              @      1@      @      1@      �?      @      �?      @                      �?      ,@                       @      @      7@      @               @      7@       @      &@      �?      �?              �?      �?              �?      $@              $@      �?                      (@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ7�+hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B6         r       	          ����?X�<ݚ�?U           ��@       /       
             �?6n�
$)�?6           `}@              	          833�?�'�`d�?g            �d@                          �b@85�}C�?L            �^@                          ``@ r���?:            �W@������������������������       �        ,             R@                           �?���}<S�?             7@       	                    �?�r����?             .@������������������������       �                     $@
                           �J@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @                           �?l��
I��?             ;@������������������������       �                     $@                          0e@��.k���?             1@                           �?�<ݚ�?             "@������������������������       �                     @              
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �?      �?              @                          �f@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                             L@�K��&�?            �E@                           _@�����H�?             2@                          �^@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     &@!       .                    �?��H�}�?             9@"       )                   �`@�\��N��?             3@#       $                   �X@�n_Y�K�?             *@������������������������       �                      @%       &                    �?���!pc�?             &@������������������������       �                     @'       (                   Pm@      �?             @������������������������       �                     @������������������������       �                     �?*       +                   `a@r�q��?             @������������������������       �                     @,       -       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @0       q                   �f@Xny��?�            s@1       B                   �O@L:�f@�?�            �r@2       9                    �?�G��l��?             5@3       4                    �?�q�q�?             "@������������������������       �                     �?5       8                   �]@      �?              @6       7                   `V@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @:       A                    �P@�q�q�?             (@;       @                    �?z�G�z�?             $@<       =                   @`@�����H�?             "@������������������������       �                     @>       ?       	          hff�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @C       P                    \@����8y�?�            �q@D       O                    �?Jm_!'1�?            �H@E       H                   Pl@     ��?             0@F       G                   �c@����X�?             @������������������������       �                     @������������������������       �                      @I       N                    �?�<ݚ�?             "@J       K                   @n@      �?              @������������������������       �                     @L       M                   �p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                    �@@Q       f                    �?�a�� �?�             m@R       e                    �?��Hg���?$            �F@S       b                    b@�(�Tw��?            �C@T       Y                    `@     ��?             @@U       V                     B@      �?              @������������������������       �                     �?W       X                    _@����X�?             @������������������������       �                     @������������������������       �                      @Z       [                   �c@�8��8��?             8@������������������������       �                     2@\       a                   0e@�q�q�?             @]       ^                    �?�q�q�?             @������������������������       �                     �?_       `                     M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @c       d                   �s@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @g       j                   `_@��p�b��?|            `g@h       i                    @P���Q�?             4@������������������������       �                     3@������������������������       �                     �?k       l                   �`@�E��La�?m            �d@������������������������       �        @             Y@m       p                    a@�\=lf�?-            �P@n       o                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        +            @P@������������������������       �                     @s       �                    �?������?            |@t       �                    �?�]z�}�?�            �r@u       �       
             �?ox%�:�?.            @R@v       �                   �a@j�q����?             I@w       �                    �N@¦	^_�?             ?@x              	          ����?�S����?             3@y       ~                    ]@      �?              @z       }       	          ����?���Q��?             @{       |                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     &@�       �                   `v@      �?             (@�       �                    �?���Q��?             $@������������������������       �                     @�       �                   @\@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     3@�       �                   pb@
;&����?             7@�       �       	          033�?     ��?             0@�       �                     L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   `T@�C��2(�?             &@������������������������       �                     "@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?���
���?�             l@�       �                    Z@�˫���?u             g@�       �                    �?r�q��?             @�       �                   �Y@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          `ff @�x�E~�?q            @f@�       �                    `R@��.N"Ҭ?T            @a@�       �                   pl@`Y����?S             a@�       �                   `_@���N8�?)            �O@������������������������       �                     E@�       �                     L@؇���X�?             5@�       �                   pb@�X�<ݺ?             2@������������������������       �                     *@�       �       	             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �i@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        *            �R@������������������������       �                     �?������������������������       �                     D@�       �                   j@��p\�?            �D@�       �                    c@z�G�z�?
             $@�       �                    �?�����H�?	             "@�       �                   �`@z�G�z�?             @�       �       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    @G@�g�y��?             ?@�       �                    ^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     =@�       �                    �?�EH,���?]            �b@�       �       
             �?և���X�?H            �]@�       �                    �D@j���� �?3            @U@������������������������       �                     @�       �                    @t�C�#��?0            �S@�       �                    �?4�	~���?)            @Q@�       �       	             �?�z�G��?             4@�       �       	          ����?؇���X�?             @�       �                    b@z�G�z�?             @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     *@�       �                    �Q@ZՏ�m|�?            �H@�       �       
             �?���H��?             E@�       �                   �_@r�q��?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�����H�?             B@������������������������       �                     @�       �                   �`@      �?             @@������������������������       �                     .@�       �                   �d@������?             1@�       �       	          ����?     ��?
             0@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �       	          `ff�?$�q-�?             *@�       �                    @M@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?�       �       	          hff@և���X�?             @�       �                    [@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @J@�z�G��?             $@������������������������       �                      @�       �                     N@      �?              @������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �]@г�wY;�?             A@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     =@�       �                   Pb@�n`���?             ?@������������������������       �                     7@�       �                   Pe@      �?              @������������������������       �                     @�       �                   @b@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp       �y@     �@     s@     �d@     �A@     @`@      $@      \@       @     @W@              R@       @      5@       @      *@              $@       @      @       @                      @               @       @      3@              $@       @      "@      @       @      @              �?       @      �?                       @      �?      @      �?       @               @      �?                      @      9@      2@      0@       @      @       @      @                       @      &@              "@      0@      "@      $@       @      @               @       @      @      @              �?      @              @      �?              �?      @              @      �?      �?              �?      �?                      @     �p@     �A@     �p@      @@      &@      $@      @      @      �?               @      @       @      �?              �?       @                      @       @      @       @       @       @      �?      @               @      �?       @                      �?              �?               @     0p@      6@      D@      "@      @      "@      @       @      @                       @       @      @      �?      @              @      �?       @      �?                       @      �?             �@@             `k@      *@      A@      &@      <@      &@      ;@      @      @      @              �?      @       @      @                       @      6@       @      2@              @       @      �?       @              �?      �?      �?      �?                      �?      @              �?      @              @      �?              @              g@       @      3@      �?      3@                      �?     �d@      �?      Y@             �P@      �?      �?      �?              �?      �?             @P@                      @     �Y@     �u@      =@     �p@      5@      J@      "@     �D@      "@      6@      @      0@      @      @      @       @      �?       @      �?                       @       @                      @              &@      @      @      @      @              @      @       @               @      @               @                      3@      (@      &@      @      &@      @      �?      @                      �?      �?      $@              "@      �?      �?      �?                      �?      @               @      k@      @     `f@      �?      @      �?       @               @      �?                      @      @     �e@      @     �`@      @     �`@      @      N@              E@      @      2@      �?      1@              *@      �?      @      �?                      @       @      �?       @                      �?             �R@      �?                      D@      @      C@       @       @      �?       @      �?      @      �?      �?      �?                      �?              @              @      �?              �?      >@      �?      �?      �?                      �?              =@     �R@      S@      Q@     �I@     �A@      I@      @              =@      I@      6@     �G@      ,@      @      �?      @      �?      @      �?      �?              �?      �?                      @               @      *@               @     �D@      @     �B@      �?      @              @      �?      �?      �?                      �?      @      @@              @      @      <@              .@      @      *@      @      *@       @      �?              �?       @              �?      (@      �?      @              @      �?                      "@      �?              @      @      @      �?              �?      @                      @      @      @               @      @      �?      @              �?      �?              �?      �?             �@@      �?      @      �?              �?      @              =@              @      9@              7@      @       @      @              �?       @               @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��mohG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B(<         �                   pb@n�A��?N           ��@       [                    �?���-���?f           `�@                          `\@X�̔���?�            �q@                           @E@v���EO�?-            �Q@������������������������       �                     @                           �?�z����?+            @P@                          �\@��}*_��?             ;@������������������������       �                      @	       
                    �?`�Q��?             9@������������������������       �                     �?              
             �?�q�q�?             8@                           �?      �?             0@������������������������       �        
             .@������������������������       �                     �?                           X@      �?              @������������������������       �                     �?������������������������       �                     @              
             �?P�Lt�<�?             C@������������������������       �                     A@              	          ����?      �?             @������������������������       �                     @������������������������       �                     �?       2                    �?r���@�?�            �j@       )       
             �?���y�?8            @V@       (                    �?"pc�
�?$            �K@                           �?�E��ӭ�?             B@                          �a@���|���?             &@������������������������       �                     @������������������������       �                     @                            O@H%u��?             9@������������������������       �                     ,@        !       	             �?���!pc�?             &@������������������������       �                     @"       '                     P@և���X�?             @#       $       	          `ff�?      �?             @������������������������       �                     �?%       &       
             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@*       -                   �`@ҳ�wY;�?             A@+       ,                    P@     ��?             0@������������������������       �                     @������������������������       �                     *@.       1       	          hff�?      �?             2@/       0                   @E@"pc�
�?             &@������������������������       �                      @������������������������       �                     "@������������������������       �                     @3       P                    �P@z�G�z�?L            @_@4       E                    @�`�=	�?A            �Y@5       @                   �_@t��ճC�?6             V@6       7                   `_@�Ra����?             F@������������������������       �                     ,@8       ;       
             �?r�q��?             >@9       :                   �a@���Q��?             @������������������������       �                     @������������������������       �                      @<       =       	          @33�?HP�s��?             9@������������������������       �                     6@>       ?                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?A       B                    �L@`���i��?             F@������������������������       �                     >@C       D                   Pj@@4և���?             ,@������������������������       �                     *@������������������������       �                     �?F       G       
             �?��S���?             .@������������������������       �                     @H       O                    �?�q�q�?	             (@I       J                    �?      �?              @������������������������       �                     @K       L                   �`@z�G�z�?             @������������������������       �                      @M       N                    a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @Q       X                    �?      �?             6@R       W                    @z�G�z�?             $@S       T                    �?�����H�?             "@������������������������       �                     @U       V       	          hff@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?Y       Z                    �R@      �?             (@������������������������       �                     "@������������������������       �                     @\       u                   i@XF�����?�            �p@]       t                    �?P���Q�?D             Y@^       s                    �?`-�I�w�?6             S@_       j       
             �?0��_��?#            �J@`       a       	          033�?�nkK�?             G@������������������������       �                     4@b       c                   �U@$�q-�?             :@������������������������       �                     �?d       e                    �?`2U0*��?             9@������������������������       �                     @f       g                   @e@P���Q�?             4@������������������������       �                     ,@h       i       	             �?r�q��?             @������������������������       �                     �?������������������������       �                     @k       l                   �Z@և���X�?             @������������������������       �                      @m       n                    �I@���Q��?             @������������������������       �                     �?o       p                    �?      �?             @������������������������       �                     �?q       r                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     7@������������������������       �                     8@v       �       	          033�?��Sa+��?q            `e@w       |                   �j@��Sݭg�?5            �S@x       y       	             �?�z�G��?             $@������������������������       �                      @z       {                   �i@      �?              @������������������������       �                     �?������������������������       �                     @}       ~                    @D@�����?/             Q@������������������������       �                     �?       �       
             �?�Y����?.            �P@�       �                    �?      �?'             L@������������������������       �                     ,@�       �                    @K@r�q��?             E@������������������������       �                     2@�       �       	          ����?�q�q�?             8@�       �       	             �?j���� �?             1@������������������������       �                     @�       �                   �q@��
ц��?	             *@�       �                   0p@      �?              @�       �                   @`@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       	          ����?�eP*L��?             &@������������������������       �                     @�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �       	          ���@�g�y��?<            @W@�       �                   0i@`����֜?,            �Q@������������������������       �                     �?������������������������       �        +            @Q@�       �                    �?���}<S�?             7@������������������������       �        
             ,@�       �                   �`@�<ݚ�?             "@�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?8�{�?�            �v@�       �                   Pe@�n\�GZ�?H            �]@�       �                    T@�����?<            �W@������������������������       �                     ,@�       �                   �b@��}*_��?4            @T@�       �                    �M@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�       �                    �?�z�G��?0            �Q@�       �       	             @:���W�?)            �M@�       �                   �i@j���� �?$            �I@�       �                   �b@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?      �?             D@�       �                    d@ҳ�wY;�?
             1@�       �                    �?�q�q�?             "@�       �                   y@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                   �r@�û��|�?             7@�       �                    `@��.k���?             1@�       �                     N@"pc�
�?
             &@�       �                   pj@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     &@�       �                    �?�q�q�?             8@�       �                    �D@8����?             7@�       �                   �f@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?���y4F�?	             3@�       �       	          @33�?r�q��?             2@�       �                   0f@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     "@������������������������       �                     �?������������������������       �                     �?�       �                   �O@T$�#���?�            `n@�       �       	            �?�eP*L��?             &@������������������������       �                     @�       �                    �N@����X�?             @������������������������       �                     @������������������������       �                      @�       �       
             �?\-��p�?�             m@�       �       
             �?T�7�s��?,            �L@������������������������       �                     @�       �                   �_@��B����?'             J@�       �                    �?`�Q��?             9@�       �                   �]@�GN�z�?             6@�       �       	          @33�?ףp=
�?             $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �n@�q�q�?             (@������������������������       �                     @�       �                    �?z�G�z�?             @�       �                    �K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	          ����?��}*_��?             ;@�       �       	          ����?�eP*L��?             6@�       �                   pc@p�ݯ��?             3@�       �                    @N@r�q��?             @�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   ``@8�Z$���?	             *@������������������������       �                     �?�       �                    �?�8��8��?             (@�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�                         �s@`2U0*��?n            �e@                          @L@PL��V�?`            �b@������������������������       �        O             _@      	                   c@      �?             8@            	            �?�}�+r��?             3@������������������������       �        
             .@                         �O@      �?             @                        @g@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @
                        Pc@���Q��?             @������������������������       �                      @������������������������       �                     @                         @L@PN��T'�?             ;@������������������������       �        	             2@            	          ����?X�<ݚ�?             "@                         `@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KMKK��h_�B0       �z@     �~@      f@     �w@     �b@      a@      1@      K@      @              &@      K@      $@      1@       @               @      1@              �?       @      0@      �?      .@              .@      �?              @      �?              �?      @              �?     �B@              A@      �?      @              @      �?             �`@     �T@      @@     �L@      $@     �F@      $@      :@      @      @      @                      @      @      6@              ,@      @       @              @      @      @      @      @      �?               @      @       @                      @              �?              3@      6@      (@      *@      @              @      *@              "@      "@      "@       @               @      "@                      @      Y@      9@     @V@      ,@     �T@      @     �C@      @      ,@              9@      @       @      @              @       @              7@       @      6@              �?       @               @      �?             �E@      �?      >@              *@      �?      *@                      �?      @       @      @              @       @      @      @      @              �?      @               @      �?       @               @      �?                      @      &@      &@       @       @       @      �?      @              @      �?      @                      �?              �?      @      "@              "@      @              <@     `n@      @     �W@      @     �Q@      @      H@       @      F@              4@       @      8@      �?              �?      8@              @      �?      3@              ,@      �?      @      �?                      @      @      @               @      @       @              �?      @      �?      �?               @      �?       @                      �?              7@              8@      7@     �b@      4@      M@      @      @               @      @      �?              �?      @              *@     �K@      �?              (@     �K@      @     �H@              ,@      @     �A@              2@      @      1@      @      $@              @      @      @      @      @      @      �?              �?      @                      @      @      �?      �?      �?              �?      �?              @                      @      @      @      @              �?      @              @      �?              @     �V@      �?     @Q@      �?                     @Q@       @      5@              ,@       @      @       @      �?       @                      �?              @     �o@     �[@      G@     @R@      >@     @P@              ,@      >@     �I@      "@       @      "@                       @      5@     �H@      5@      C@      5@      >@      �?      $@              $@      �?              4@      4@      @      &@      @      @      @      �?      @                      �?       @       @       @                       @               @      ,@      "@       @      "@       @      "@      �?       @      �?                       @      �?      �?              �?      �?              @              @                       @              &@      0@       @      0@      @      �?      @              @      �?              .@      @      .@      @      @      @              @      @              "@                      �?              �?     �i@     �B@      @      @      @               @      @              @       @              i@      @@      @@      9@      @              ;@      9@      1@       @      1@      @      "@      �?      �?      �?      �?                      �?       @               @      @      @              �?      @      �?       @      �?                       @               @              @      $@      1@      $@      (@      @      (@      @      �?      �?      �?      �?                      �?      @               @      &@      �?              �?      &@      �?      @      �?                      @              @      @                      @      e@      @      b@      @      _@              5@      @      2@      �?      .@              @      �?      �?      �?      �?                      �?       @              @       @               @      @              7@      @      2@              @      @      �?      @      �?                      @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ2LAVhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�:         �                    �?Ь�g���?;           ��@                          @E@JZ�]�[�?4           0~@                          �V@��(\���?L             ^@������������������������       �                      @                          �Z@�1e�3��?K            �]@������������������������       �                    �@@                          �Z@�m(�X�?3            @U@������������������������       �                     �?	                           �?@4և���?2             U@
                           �?�<ݚ�?             ;@                          p`@�����H�?             2@������������������������       �        
             .@                           �?�q�q�?             @������������������������       �                     �?������������������������       �                      @              
             �?X�<ݚ�?             "@              
             �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @                           �I@      �?             @                            E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                    �L@       M                    �?����ƛ�?�            �v@       (                   P`@^�tD|��?V            �a@       !                    �?r�z-��?!            �J@                           �E@r�q��?             (@������������������������       �                     �?                           �`@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?"       '       	             �?� ��1�?            �D@#       &       
             �?������?             >@$       %                    U@�nkK�?             7@������������������������       �                     �?������������������������       �                     6@������������������������       �                     @������������������������       �        	             &@)       H                   �s@�μ���?5            @V@*       +                   pd@̘SJl��?0            �S@������������������������       �                     $@,       G       	          ���@��<b���?,            @Q@-       0                    �?�'݊U�?*            �P@.       /                   �b@���N8�?             5@������������������������       �        
             4@������������������������       �                     �?1       :                    �?��+7��?             G@2       3                    @F@�eP*L��?             &@������������������������       �                      @4       5                   �j@�q�q�?             "@������������������������       �                     �?6       7                   �a@      �?              @������������������������       �                     @8       9                    ^@���Q��?             @������������������������       �                     @������������������������       �                      @;       F                   �l@z�G�z�?            �A@<       E                    @J@p�ݯ��?             3@=       >                   �b@��
ц��?	             *@������������������������       �                     @?       @                   0k@�z�G��?             $@������������������������       �                     @A       D                   �l@      �?             @B       C                   @b@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     0@������������������������       �                      @I       J                    �E@�z�G��?             $@������������������������       �                      @K       L                    �?      �?              @������������������������       �                     �?������������������������       �                     @N       s       	          ����?�K�̀��?�            �k@O       r                    �?�q�q�?/             R@P       o                   �s@�z�G��?$             I@Q       n                   �r@��+7��?!             G@R       Y                   @\@�q�q�?             B@S       T                    �I@���Q��?             $@������������������������       �                      @U       V                    k@      �?              @������������������������       �                     �?W       X       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?Z       c                    �?�θ�?             :@[       `       	          433�?�q�q�?             "@\       ]                   @n@      �?             @������������������������       �                      @^       _                   �n@      �?              @������������������������       �                     �?������������������������       �                     �?a       b                    a@���Q��?             @������������������������       �                      @������������������������       �                     @d       i                   �`@@�0�!��?             1@e       f                     N@ףp=
�?	             $@������������������������       �                      @g       h       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?j       m                    �G@����X�?             @k       l                    @D@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     $@p       q       
             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     6@t       w                   �Z@ཕvt�?c            �b@u       v                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?x       �                   pb@@9G��?a            `b@y       �                    _@ T���v�?I            @\@z       �                   pp@      �?             @@{       �                   �o@�����?             5@|       }       
             �?P���Q�?             4@������������������������       �                     @~       �       	          ����?�IєX�?             1@       �                     M@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@������������������������       �                     �?������������������������       �                     &@�       �                   �b@ �)���?3            @T@������������������������       �        .            �Q@�       �                    q@�C��2(�?             &@������������������������       �                     @�       �                   �q@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �       	             @l��\��?             A@�       �                    �R@     ��?
             0@�       �                   �_@@4և���?	             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                      @������������������������       �                     2@�       �                    �?������?           0{@�       �                   �c@��!����?�            �v@�       �       
             �?8����?             G@�       �                    `Q@�חF�P�?             ?@�       �                    �?@4և���?             <@������������������������       �                     �?�       �                   �Q@ 7���B�?             ;@������������������������       �                     4@�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       	            �?���Q��?             .@�       �                     Q@"pc�
�?             &@������������������������       �                      @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?R���Q�?�             t@�       �                    �?L��B�?�            �q@�       �                   r@������?!             K@�       �                    @L@�q�q�?             H@�       �                   pg@XB���?             =@������������������������       �                     <@������������������������       �                     �?�       �       	          033�?�����?             3@�       �                    q@��
ц��?             *@�       �                    @M@���Q��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       
             �?�J��?�            �l@�       �       	          `ff�?     ��?             @@�       �                   �Z@�+e�X�?             9@������������������������       �                     �?�       �       	          ����?�q�q�?             8@�       �                    @�t����?             1@�       �                    �?      �?             0@�       �                   0q@�C��2(�?	             &@������������������������       �                     $@������������������������       �                     �?�       �                    j@���Q��?             @������������������������       �                     �?�       �                     K@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �`@����X�?             @�       �                   @_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �O@���p�T�?v            �h@�       �                    @L@@�Ջ��?q            �g@�       �                   @[@�����?e            �e@�       �                    �G@$�q-�?             *@�       �                   �c@      �?             @�       �                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �        ^             d@�       �                    �?�����H�?             2@������������������������       �                      @�       �       	            �?z�G�z�?             $@������������������������       �                     @�       �                   a@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �s@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                     H@��+��?            �B@������������������������       �                     "@�       �                    �?X�Cc�?             <@�       �                   �[@�G��l��?             5@������������������������       �                      @�       �                    @D�n�3�?             3@�       �                   0k@b�2�tk�?             2@������������������������       �                      @�       �       	             �?     ��?
             0@�       �                   �\@�q�q�?             (@������������������������       �                      @�       �       
             �?�z�G��?             $@�       �                   �r@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�                          �?
;&����?*            @Q@�                         �c@���Q��?             I@�       �                   �`@�X����?             F@������������������������       �                     @�       �       	            �?���� �?            �D@�       �       
             �?PN��T'�?             ;@������������������������       �                     @������������������������       �                     7@�       �                    @L@      �?
             ,@������������������������       �                     @�              
             �?���|���?             &@������������������������       �                     @                         �?z�G�z�?             @������������������������       �                     @                         �M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        Pj@�S����?             3@������������������������       �                     &@	                         �?      �?              @
                        �o@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�t�b�j"     h�h(h+K ��h-��R�(KMKK��h_�B�       0{@     0~@      ]@     �v@      "@     �[@       @              @     �[@             �@@      @     �S@      �?              @     �S@      @      5@       @      0@              .@       @      �?              �?       @              @      @      �?      @      �?                      @      @      �?      �?      �?      �?                      �?       @                     �L@     �Z@      p@     @U@     �L@      2@     �A@      $@       @              �?      $@      �?      $@                      �?       @     �@@       @      6@      �?      6@      �?                      6@      @                      &@     �P@      6@      P@      .@      $@              K@      .@      K@      *@      4@      �?      4@                      �?      A@      (@      @      @               @      @      @              �?      @       @      @              @       @      @                       @      <@      @      (@      @      @      @      @              @      @              @      @      @      @      �?      @                      �?               @      @              0@                       @      @      @       @              �?      @      �?                      @      6@     �h@      .@     �L@      .@     �A@      (@      A@      (@      8@      @      @               @      @       @              �?      @      �?      @                      �?      @      4@      @      @      �?      @               @      �?      �?      �?                      �?       @      @       @                      @      @      ,@      �?      "@               @      �?      �?      �?                      �?       @      @       @      �?              �?       @                      @              $@      @      �?      @                      �?              6@      @     �a@      �?      �?              �?      �?              @     �a@      @     �[@       @      >@       @      3@      �?      3@              @      �?      0@      �?      @      �?                      @              (@      �?                      &@      �?      T@             �Q@      �?      $@              @      �?      @      �?                      @      @      ?@      @      *@      �?      *@              *@      �?               @                      2@     �s@      ]@     �q@      T@      ,@      @@      @      :@       @      :@      �?              �?      :@              4@      �?      @      �?                      @      @              "@      @      "@       @       @              �?       @      �?                       @              @      q@      H@     �o@      >@      D@      ,@      A@      ,@      <@      �?      <@                      �?      @      *@      @      @      @      @              @      @                      @              @      @             �j@      0@      5@      &@      3@      @              �?      3@      @      (@      @      (@      @      $@      �?      $@                      �?       @      @      �?              �?      @              �?      �?       @      �?                       @              �?      @               @      @       @       @               @       @                      @      h@      @     �g@      @     �e@      �?      (@      �?      @      �?      �?      �?      �?                      �?       @              "@              d@              0@       @       @               @       @      @               @       @               @       @              @       @      @                       @      3@      2@      "@              $@      2@      $@      &@       @               @      &@      @      &@               @      @      "@      @      @               @      @      @      @      @              @      @              @                      @      �?                      @     �@@      B@      >@      4@      >@      ,@              @      >@      &@      7@      @              @      7@              @      @      @              @      @              @      @      �?      @              �?      �?      �?                      �?              @      @      0@              &@      @      @      @      �?      @                      �?              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJو�1hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�Bx=         �       
             �?z�ГPo�?T           ��@       y                   �b@��8Y.��?N           �@       <                    �?��]�?           0z@                          `\@�<ݚ�?T            �_@                          `x@`Ӹ����?            �F@                           �?`���i��?             F@                          @^@�nkK�?             7@       	                    �K@؇���X�?             @������������������������       �                     @
                          �X@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        	             0@������������������������       �                     5@������������������������       �                     �?       ;                    �?�w���?7            @T@       "                    @J@lutee�?+            �P@                          �f@"pc�
�?            �@@������������������������       �                     @                           �?�θ�?             :@                           @H@�KM�]�?	             3@������������������������       �                     &@              	             �?      �?              @������������������������       �                     @                          �`@      �?             @������������������������       �                      @������������������������       �                      @                           k@և���X�?             @������������������������       �                     @       !                   @b@      �?             @                            �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @#       :                   @q@j���� �?             A@$       '                    [@      �?             @@%       &                   �f@      �?             @������������������������       �                     @������������������������       �                     �?(       )       	          ����?��X��?             <@������������������������       �                     @*       /                   �k@�q�q�?             8@+       ,                   pj@��S�ۿ?	             .@������������������������       �                     $@-       .                    k@z�G�z�?             @������������������������       �                     �?������������������������       �                     @0       1       	          hff�?X�<ݚ�?             "@������������������������       �                     �?2       3       
             �?      �?              @������������������������       �                     �?4       5                   0b@և���X�?             @������������������������       �                     @6       7                    �?      �?             @������������������������       �                      @8       9                   Pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@=       P                    �?�yI�n�?�            Pr@>       O                    �?д>��C�?             =@?       B       	          ����?z�G�z�?             9@@       A                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @C       D                    �?��2(&�?             6@������������������������       �                     @E       N                   �r@@�0�!��?             1@F       M       	          ����?���!pc�?	             &@G       L                    �?և���X�?             @H       K                   �m@�q�q�?             @I       J                     M@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @Q       v                   `f@ �q�q�?�            �p@R       i                    �?����?�            @p@S       \                    �? _�@�Y�?�             m@T       U                   �_@@�����?g             e@������������������������       �        C            @\@V       [       	          ����?�h����?$             L@W       X       	          ����?���7�?             6@������������������������       �                     4@Y       Z                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     A@]       b                   �_@���N8�?)            �O@^       _       	             @�<ݚ�?             "@������������������������       �                     @`       a                   �^@���Q��?             @������������������������       �                     @������������������������       �                      @c       h                    �L@@3����?%             K@d       g                   �Z@ �q�q�?             8@e       f                    b@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     3@������������������������       �                     >@j       o                   �[@�>4և��?             <@k       l                    �?���Q��?             @������������������������       �                     �?m       n                   �Z@      �?             @������������������������       �                      @������������������������       �                      @p       u       	          ����?���}<S�?             7@q       r                   �l@z�G�z�?             $@������������������������       �                     @s       t                   @[@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@w       x                   �X@      �?             @������������������������       �                      @������������������������       �                      @z       �                    �?֦�r��?<            �U@{       �                    �?$�q-�?            �C@|                          pc@R���Q�?             4@}       ~       	             @�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �e@�IєX�?
             1@������������������������       �        	             0@������������������������       �                     �?������������������������       �                     3@�       �                    �?(���@��?#            �G@�       �                   `a@\�Uo��?             C@�       �                   `l@8^s]e�?             =@�       �                    �L@@4և���?
             ,@������������������������       �                     &@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?��S���?             .@�       �                   0f@      �?             ,@�       �                    e@�z�G��?             $@�       �                    @K@և���X�?             @������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                     O@�q�q�?             "@�       �                   f@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@�       �                    �L@x�͛��?           �y@�       �       	            �?�Qb��?�            �r@�       �                    �?���C���?�             o@�       �                   @E@     ��?%             P@�       �                    �J@      �?              @�       �                    @I@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                    �?�>4և��?!             L@�       �                   �c@��Q��?             4@�       �                    n@�eP*L��?             &@�       �                     G@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    ]@�����H�?             "@�       �                    e@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   pf@�8��8��?             B@�       �                    `@г�wY;�?             A@�       �                   �o@$�q-�?             *@������������������������       �                      @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     5@������������������������       �                      @�       �                    �?hl �&�?z             g@�       �                   �g@H%u��?             9@������������������������       �                     4@�       �                    �D@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   @n@�O4R���?j            �c@������������������������       �        @            �X@�       �                   �n@P���Q�?*             N@������������������������       �                     @������������������������       �        )            �L@�       �                    `@�>���?"             K@�       �                   @^@      �?             @@�       �                   �f@�G��l��?             5@������������������������       �                      @�       �                    b@8�Z$���?             *@�       �                   �o@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @�       �                    �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �                    �?�GN�z�?             6@�       �                   �V@      �?             $@������������������������       �                      @�       �                   Pc@      �?              @�       �                    �?      �?             @������������������������       �                      @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       �                   �]@��J�fj�?E            �[@�       �                   �[@���N8�?             5@�       �       	          ����?�eP*L��?             &@�       �                   @Y@����X�?             @�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     $@�             	          ����?�L�lRT�?9            �V@�                         �f@�d�����?0             S@�       �                    �?���"͏�?/            �R@�       �                    �?d��0u��?             >@�       �                    b@R�}e�.�?             :@�       �                    �?؇���X�?             ,@������������������������       �                     $@�       �                   0`@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �\@�q�q�?             (@������������������������       �                     @�       �                   `Y@�<ݚ�?             "@������������������������       �                     @�       �                   �c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�                          �O@fP*L��?             F@�                         `c@ܷ��?��?             =@�       �                   @b@$�q-�?             :@������������������������       �                     &@�                           �?�r����?	             .@�       �                   @a@r�q��?             (@������������������������       �                      @������������������������       �                     $@������������������������       �                     @                         �?�q�q�?             @������������������������       �                      @������������������������       �                     �?      
                  �c@������?             .@                         �Q@�C��2(�?	             &@������������������������       �                      @      	                   `R@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         d@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @                        @l@؇���X�?	             ,@                         @N@�8��8��?             (@                         �?      �?             @                        �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                        p`@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KMKK��h_�B�       �x@     @�@     �S@     �z@      F@     pw@      <@     �X@       @     �E@      �?     �E@      �?      6@      �?      @              @      �?      @      �?                      @              0@              5@      �?              :@     �K@      :@     �D@      @      ;@              @      @      4@       @      1@              &@       @      @              @       @       @       @                       @      @      @      @              �?      @      �?      �?      �?                      �?               @      4@      ,@      4@      (@      �?      @              @      �?              3@      "@              @      3@      @      ,@      �?      $@              @      �?              �?      @              @      @      �?              @      @      �?              @      @              @      @      �?       @              �?      �?      �?                      �?               @              ,@      0@     Pq@      @      8@      @      4@       @      �?              �?       @              @      3@              @      @      ,@      @       @      @      @       @      @       @      �?       @                      �?              @      �?                      @              @              @      &@     �o@      "@     `o@      @     �l@      �?      e@             @\@      �?     �K@      �?      5@              4@      �?      �?              �?      �?                      A@      @      N@       @      @              @       @      @              @       @              �?     �J@      �?      7@      �?      @      �?                      @              3@              >@      @      7@      @       @      �?               @       @               @       @               @      5@       @       @              @       @      �?              �?       @                      *@       @       @       @                       @     �A@     �I@      @      B@      @      1@       @      �?       @                      �?      �?      0@              0@      �?                      3@      @@      .@      7@      .@      4@      "@      *@      �?      &@               @      �?              �?       @              @       @      @      @      @      @      @      @       @              �?      @      �?                      @              @      @                      �?      @      @      �?      @              @      �?               @              "@             �s@     �W@      p@      G@     `l@      5@     �H@      .@      @      @      @       @               @      @                      @      G@      $@      *@      @      @      @      @      �?              �?      @                      @       @      �?       @      �?       @                      �?      @             �@@      @     �@@      �?      (@      �?       @              @      �?      @                      �?      5@                       @     @f@      @      6@      @      4@               @      @       @                      @     �c@      @     �X@             �L@      @              @     �L@              =@      9@      (@      4@      &@      $@               @      &@       @      @       @               @      @               @              �?      $@              $@      �?              1@      @      @      @               @      @      @      �?      @               @      �?      �?      �?                      �?      @              (@             �O@      H@      @      0@      @      @      @       @      �?       @      �?                       @      @                      @              $@      M@      @@      L@      4@      L@      2@      3@      &@      3@      @      (@       @      $@               @       @       @                       @      @      @              @      @       @      @               @       @       @                       @              @     �B@      @      :@      @      8@       @      &@              *@       @      $@       @               @      $@              @               @      �?       @                      �?      &@      @      $@      �?       @               @      �?              �?       @              �?      @              @      �?                       @       @      (@      �?      &@      �?      @      �?      �?      �?                      �?               @               @      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK݅�h~�BX0         z       	          033�?>���i��?I           ��@       -       
             �?�\�J��?>           p@              	          ����?� ��1�?k            �d@                           �?`Jj��?O             _@                           �?����X�?             5@                          @a@      �?             @������������������������       �                     �?������������������������       �                     @	                          �c@@�0�!��?             1@
                           �G@@4և���?             ,@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@                           @F@�q�q�?             @������������������������       �                     �?                          8p@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?p� V�?B            �Y@������������������������       �        /             R@              
             �?`Jj��?             ?@������������������������       �                     �?                           Z@(;L]n�?             >@                          `Z@      �?              @                           X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@       "       	          ����?���Q��?             D@        !                    X@�����H�?
             2@������������������������       �                      @������������������������       �        	             0@#       $                    �?���|���?             6@������������������������       �                     @%       ,                    �?@�0�!��?             1@&       '       
             �?և���X�?             @������������������������       �                      @(       )                    �?z�G�z�?             @������������������������       �                     @*       +                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@.       ]                    �?4Ky\�?�            0u@/       R                    �?�q�q��?;             X@0       E                    �K@��cv�?/            @S@1       4                    P@r֛w���?$             O@2       3                    �?r�q��?             @������������������������       �                     @������������������������       �                     �?5       D                   0o@����>4�?!             L@6       7                   �a@<ݚ)�?             B@������������������������       �        	             1@8       C                   �f@D�n�3�?             3@9       :                    �?b�2�tk�?             2@������������������������       �                      @;       B                    �?�z�G��?             $@<       A                    @J@�q�q�?             "@=       @                   @b@      �?             @>       ?                   `l@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@F       Q                    �?��S���?             .@G       H                    i@���|���?	             &@������������������������       �                     @I       P       	          ����?      �?              @J       K                   �`@և���X�?             @������������������������       �                      @L       M                   �i@���Q��?             @������������������������       �                      @N       O                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @S       \                     O@�d�����?             3@T       U                   �Z@      �?             $@������������������������       �                     @V       Y                   �`@����X�?             @W       X                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?Z       [                    �K@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@^       q                   �s@�g�H��?�            `n@_       n                    �Q@h�����?�             l@`       e                   @[@ �� ��?�            �k@a       d                    �G@؇���X�?             ,@b       c                   �Z@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @f       g       	            �?@$��g�?�            �i@������������������������       �        o             f@h       i                   @d@�r����?             >@������������������������       �                     �?j       k                    @L@ܷ��?��?             =@������������������������       �                     3@l       m                     O@�z�G��?             $@������������������������       �                     @������������������������       �                     @o       p                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @r       y                    d@�d�����?             3@s       t                    @L@�n_Y�K�?             *@������������������������       �                     @u       x                    �?����X�?             @v       w                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @{       �                    �?�� ���?           �y@|       �                   �g@X9����?V            �_@}       ~                   `_@��E�B��?#            �G@������������������������       �                     1@       �                   �c@z�G�z�?             >@�       �                    �?ȵHPS!�?             :@�       �                    T@�z�G��?             $@�       �       	          hff@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     0@�       �                    `@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?��Q���?3             T@�       �       	             �?���@M^�?             ?@�       �                   �l@ҳ�wY;�?	             1@������������������������       �                     @������������������������       �                     &@�       �                    n@@4և���?	             ,@�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �       	          ���@ZՏ�m|�?!            �H@�       �       	             �?��p\�?            �D@�       �       
             �?     ��?	             0@�       �                   Xs@      �?             @�       �       	          ����?      �?             @������������������������       �                      @�       �       	          pff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     9@�       �                    �?      �?              @������������������������       �                     �?�       �       	             
@����X�?             @������������������������       �                     @�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @�����H�?�             r@�       �                   P`@�d�g��?�            �q@�       �                   �h@�חF�P�?O             _@������������������������       �                     B@�       �                   �m@�GN�z�?6             V@�       �                   `a@؀�:M�?            �B@�       �                   �\@��2(&�?             6@�       �                    �I@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   @X@�}�+r��?             3@������������������������       �                     �?������������������������       �                     2@�       �                    �?������?             .@������������������������       �                     &@������������������������       �                     @�       �                    �?�t����?            �I@�       �                   ``@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                   �\@����?�?            �F@�       �                    �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                    �@@�       �                    �? ��WV�?a            �c@�       �                   pl@z�G�z�?             .@�       �                   �j@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                     E@`Ql�R�?U            �a@�       �                   �g@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    c@ aqk+�?S            `a@�       �                    �?���б�?P            �`@������������������������       �        E             \@�       �                    X@�nkK�?             7@�       �                    �?�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@�       �                    �?      �?             @�       �                    �K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �a@      �?              @�       �       	          `ff@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@      t@     �f@      @@     �`@       @      ]@      @      .@      @      �?              �?      @              @      ,@      �?      *@      �?       @               @      �?                      &@       @      �?      �?              �?      �?              �?      �?               @     @Y@              R@       @      =@      �?              �?      =@      �?      @      �?       @               @      �?                      @              6@      8@      0@      0@       @               @      0@               @      ,@      @              @      ,@      @      @       @              �?      @              @      �?      �?      �?                      �?              $@      r@     �I@      M@      C@     �J@      8@      G@      0@      �?      @              @      �?             �F@      &@      9@      &@      1@               @      &@      @      &@               @      @      @      @      @      @      @      @      �?      @                      �?               @      @              �?              �?              4@              @       @      @      @      @              @      @      @      @       @               @      @               @       @      �?       @                      �?              �?              @      @      ,@      @      @              @      @       @      �?      �?      �?                      �?      @      �?      @                      �?              "@     �l@      *@      k@       @     �j@      @      (@       @      @       @      @                       @      @             `i@      @      f@              :@      @              �?      :@      @      3@              @      @              @      @              �?       @      �?                       @      ,@      @       @      @      @               @      @       @       @               @       @                      @      @             �V@     @t@     �M@      Q@      @     �D@              1@      @      8@      @      7@      @      @      @       @      @                       @              @              0@      @      �?              �?      @             �J@      ;@      (@      3@      &@      @              @      &@              �?      *@      �?      @              @      �?                      $@     �D@       @      C@      @      *@      @      @      @      �?      @               @      �?      �?      �?                      �?       @              $@              9@              @      @      �?               @      @              @       @      �?       @                      �?      @@      p@      :@     �o@      4@      Z@              B@      4@      Q@      ,@      7@      @      3@       @      �?              �?       @              �?      2@      �?                      2@      &@      @      &@                      @      @     �F@      @      �?      @                      �?      �?      F@      �?      &@              &@      �?                     �@@      @     �b@      @      (@      @      @              @      @                      "@      @     @a@      �?      �?      �?                      �?       @      a@      �?     �`@              \@      �?      6@      �?       @      �?      �?              �?      �?                      �?              4@      �?      @      �?      �?              �?      �?                       @      @       @      @      �?      @                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�6hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�6         �                    �?~jÚʞ�?8           ��@       M       
             �?��s1�?&           p~@                           �?��m�q�?�            w@                          @]@      �?!             P@������������������������       �                     (@                           `@��
ц��?             J@������������������������       �                     "@                           �J@8�$�>�?            �E@	       
       	          hff�?�	j*D�?             *@������������������������       �                     @                           �F@�q�q�?             @������������������������       �                     @                          �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?                           i@z�G�z�?             >@                          �d@�q�q�?             @������������������������       �                     @������������������������       �                      @              	          ����?�8��8��?             8@                          pc@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     .@       F                    �?�q���?�            s@                          �U@�*v��?z            @h@������������������������       �                      @       -                   @j@p�qG�?y             h@                            @L@�qM�R��?2            �P@                          �i@������?             B@������������������������       �                    �A@������������������������       �                     �?!       $                    �L@�חF�P�?             ?@"       #                   0d@      �?             @������������������������       �                     @������������������������       �                     @%       &                    �?HP�s��?             9@������������������������       �                     1@'       (                    @O@      �?              @������������������������       �                     @)       ,       
             �?���Q��?             @*       +                    X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @.       E                    �M@ ��+,��?G            @_@/       B                   0c@���N8�?1             U@0       1                    @H@x�G�z�?/             T@������������������������       �                     :@2       ;                   �\@�X�<ݺ?              K@3       :                   �a@�r����?
             .@4       9                    �?�<ݚ�?             "@5       8       	             �?      �?              @6       7                   �Y@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @<       A                    �H@ ���J��?            �C@=       @                    �?z�G�z�?             @>       ?       	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     A@C       D                   �c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                    �D@G       H                    �? �O�H�?@            �[@������������������������       �                    �C@I       L       
             �?�k~X��?'             R@J       K                   �r@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �        !             N@N       m                    �?�m����?K            �]@O       j       	             �?�E����?.             R@P       ]                    @K@�jTM��?&            �N@Q       \                   ``@<���D�?            �@@R       S       	          `ffֿ�<ݚ�?             2@������������������������       �                      @T       U                    �?      �?             0@������������������������       �                     @V       [                    �?r�q��?             (@W       X                   �b@"pc�
�?
             &@������������������������       �                     @Y       Z                   �i@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@^       i                    �?��>4և�?             <@_       f                    �?�GN�z�?             6@`       c                   �q@�S����?             3@a       b                   �a@      �?             0@������������������������       �                     .@������������������������       �                     �?d       e                    d@�q�q�?             @������������������������       �                     �?������������������������       �                      @g       h       	          @33�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @k       l                   pb@���!pc�?             &@������������������������       �                      @������������������������       �                     @n                          �q@�3Ea�$�?             G@o       t                    �I@      �?             B@p       q                    �F@����X�?             @������������������������       �                     �?r       s                   �`@r�q��?             @������������������������       �                     �?������������������������       �                     @u       ~                    @N@\-��p�?             =@v       }                   �d@��s����?             5@w       x                    �?R���Q�?             4@������������������������       �        	             &@y       z       	          `ff�?�q�q�?             "@������������������������       �                      @{       |                     M@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �       	          pff�?��� �P�?           �z@�       �       
             �?^B�z��?�             u@�       �                   �Q@t���D�?7            �U@�       �       
             �?�}�+r��?             3@������������������������       �                     �?������������������������       �                     2@�       �                   pd@B�
k���?+            �P@�       �                   hq@f�Sc��?            �H@�       �       	          ����?`՟�G��?             ?@�       �                    �K@�q�q�?             2@�       �                    �?և���X�?             @�       �                   �\@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �a@"pc�
�?             &@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                      @�       �                   �j@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �f@8�Z$���?             *@������������������������       �                     �?�       �                    @J@�8��8��?             (@�       �                    �F@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                   �X@�X�<ݺ?
             2@�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     0@�       �                   �o@�<ݚ�?             2@�       �                    �?�r����?             .@�       �                   �e@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     $@�       �                    @E@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?�i�y�?�            �o@�       �                   �d@6YE�t�?            �@@�       �                   pc@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?ףp=
�?             >@�       �                    @@4և���?             <@�       �                   pd@ ��WV�?             :@������������������������       �        
             .@�       �                   0m@�C��2(�?             &@�       �                    @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                   pl@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     R@ �й���?�            `k@�       �       	          ����?��wڝ�?�            @k@�       �                   pa@�ۘ�E-�?|            @i@������������������������       �        `            @b@�       �                    �O@�h����?             L@������������������������       �                     J@�       �                   �b@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �_@      �?
             0@������������������������       �                     �?������������������������       �        	             .@������������������������       �                     �?�       �       	          033�?4E���?>            @W@�       �                    a@�eP*L��?             F@�       �                   �_@�d�����?             3@�       �                   �\@      �?              @������������������������       �                     @�       �       	          033�?z�G�z�?             @�       �                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    Y@�C��2(�?             &@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                    �N@�+e�X�?             9@�       �                    �J@P���Q�?             4@������������������������       �                     $@�       �                   �`@ףp=
�?             $@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       
             �?�D��?"            �H@�       �                     H@      �?             @������������������������       �                      @�       �                   @]@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?>��C��?            �E@������������������������       �                     @�       �                    @F@z�G�z�?             D@�       �       	             @      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�����H�?             B@�       �       
             �?���N8�?             5@������������������������       �        
             0@�       �                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   �b@z�G�z�?
             .@������������������������       �                     "@�       �                   Pe@      �?             @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@     �W@     �x@     �B@     �t@      8@      D@              (@      8@      <@      "@              .@      <@      "@      @      @               @      @              @       @      �?       @                      �?      @      8@      @       @      @                       @       @      6@       @      @              @       @                      .@      *@     @r@      (@     �f@       @              $@     �f@      @     �N@      �?     �A@             �A@      �?              @      :@      @      @              @      @               @      7@              1@       @      @              @       @      @       @      �?       @                      �?               @      @     @^@      @      T@      @     @S@              :@      @     �I@       @      *@       @      @      �?      @      �?      �?              �?      �?                      @      �?                      @      �?      C@      �?      @      �?      @      �?                      @              �?              A@      �?      @      �?                      @             �D@      �?     �[@             �C@      �?     �Q@      �?      &@              &@      �?                      N@      M@      N@     �H@      7@      G@      .@      =@      @      ,@      @               @      ,@       @      @              $@       @      "@       @      @              @       @               @      @              �?              .@              1@      &@      1@      @      0@      @      .@      �?      .@                      �?      �?       @      �?                       @      �?       @      �?                       @              @      @       @               @      @              "@     �B@      "@      ;@      @       @              �?      @      �?              �?      @              @      9@      @      1@      @      1@              &@      @      @       @              �?      @              @      �?              �?                       @              $@     �s@     @]@     Pq@     �N@     �@@     �J@      �?      2@      �?                      2@      @@     �A@      2@      ?@      1@      ,@      @      (@      @      @      @      �?              �?      @                       @       @      "@              @       @      @               @       @      �?              �?       @              &@       @              �?      &@      �?      @      �?      @                      �?       @              �?      1@      �?      �?              �?      �?                      0@      ,@      @      *@       @      @       @               @      @              $@              �?       @      �?                       @     �n@       @      <@      @      �?       @               @      �?              ;@      @      :@       @      9@      �?      .@              $@      �?      �?      �?      �?                      �?      "@              �?      �?      �?                      �?      �?      �?              �?      �?              k@      @      k@       @      i@      �?     @b@             �K@      �?      J@              @      �?              �?      @              .@      �?              �?      .@                      �?     �B@      L@      8@      4@      @      ,@      @      @              @      @      �?       @      �?              �?       @               @              �?      $@      �?      �?              �?      �?                      "@      3@      @      3@      �?      $@              "@      �?      @      �?      @                      �?      @                      @      *@      B@      @      @       @              �?      @      �?                      @      $@     �@@      @              @     �@@      @      �?      @                      �?      @      @@      �?      4@              0@      �?      @              @      �?              @      (@              "@      @      @      @                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �                    �?<qn�h��?:           ��@       S                    @L@R��@k�?X           x�@                          `Z@�e4h�D�?�            �w@                            J@ףp=
�?             4@                           ^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     1@	       H       	          033�?����%n�?�            pv@
       #                    �?⚩ �x�?�            0t@                           �?)O���?-             R@              
             �?�q�q�?%             N@                          �^@XB���?             =@                          Pr@�IєX�?
             1@������������������������       �        	             0@������������������������       �                     �?������������������������       �                     (@                           @F@��a�n`�?             ?@                          �r@j���� �?
             1@                           �E@�q�q�?             (@                           @D@����X�?             @                           �B@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �        	             ,@                          �a@      �?             (@������������������������       �                      @                            �G@      �?             @������������������������       �                      @!       "                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?$       ;       
             �?��N*tt�?�            `o@%       &                    �?�θ�?            �C@������������������������       �        	             0@'       ,                   @b@�û��|�?             7@(       )                   �[@z�G�z�?             @������������������������       �                     @*       +                     I@      �?              @������������������������       �                     �?������������������������       �                     �?-       :                    �?�E��ӭ�?             2@.       1       	          ����?�q�q�?
             .@/       0                    @z�G�z�?             $@������������������������       �                      @������������������������       �                      @2       3       
             �?���Q��?             @������������������������       �                     �?4       7                    �?      �?             @5       6       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?8       9                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @<       ?                   `R@@䯦s#�?�            �j@=       >       	          ����?؇���X�?             @������������������������       �                     @������������������������       �                     �?@       G                   @[@����?|            �i@A       B                   �l@$�q-�?
             *@������������������������       �                      @C       D                    �?z�G�z�?             @������������������������       �                      @E       F                     H@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        r             h@I       J                    �?      �?             B@������������������������       �                     @K       L                   �d@�eP*L��?            �@@������������������������       �                      @M       R                     I@���Q��?             9@N       Q       
             �?X�<ݚ�?
             2@O       P                   �d@�θ�?             *@������������������������       �                     $@������������������������       �                     @������������������������       �                     @������������������������       �                     @T       c                   �d@��,���?s            �f@U       \                    �?���c�H�?"            �H@V       W                    @O@և���X�?             ,@������������������������       �                     @X       Y                   �`@z�G�z�?             $@������������������������       �                     @Z       [                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @]       ^                   �c@�#-���?            �A@������������������������       �                     >@_       b                    �?���Q��?             @`       a                   �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @d       �       	          ����?vA����?Q            ``@e       ~                     P@P����?.             S@f       m                   �k@>4և���?#             L@g       h                   �h@�LQ�1	�?             7@������������������������       �                     &@i       l                    �N@      �?             (@j       k                   �j@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @n       }                    b@����e��?            �@@o       |                    @O@�q�����?             9@p       {                   �`@8�A�0��?             6@q       t                   �^@     ��?
             0@r       s                    n@z�G�z�?             @������������������������       �                     �?������������������������       �                     @u       v                   �_@���!pc�?             &@������������������������       �                     @w       x       
             �?      �?              @������������������������       �                      @y       z                    �M@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @       �                   �[@R���Q�?             4@������������������������       �                     �?�       �                    j@�KM�]�?
             3@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@�       �                   �b@��N`.�?#            �K@�       �                   `v@tk~X��?             B@�       �                    �?     ��?             @@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   b@��S�ۿ?             >@�       �                    �? 7���B�?             ;@������������������������       �        	             0@�       �                   pl@�C��2(�?             &@������������������������       �                     @�       �                   0b@z�G�z�?             @������������������������       �                     @�       �       	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   0b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �c@D�n�3�?             3@�       �                    @      �?	             0@�       �                   �c@z�G�z�?             $@������������������������       �                     @�       �                   (p@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       
             �?`�5�χ�?�            pv@�       �                   �b@������?�            `s@�       �                   `_@h�Y���?�            Pr@�       �       	          `ff�?���!5��?o            `f@�       �                    �?p��@���?3            @U@�       �       	          ����? >�֕�?)            �Q@������������������������       �                     8@�       �                   �k@���}<S�?             G@������������������������       �                     7@�       �                    �?�㙢�c�?             7@������������������������       �                     @�       �                   �p@z�G�z�?             4@�       �                   �`@�q�q�?             @������������������������       �                     �?�       �                   `m@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�t����?             1@�       �                   �q@"pc�
�?             &@������������������������       �                     @�       �                   �r@����X�?             @������������������������       �                     �?�       �                   @_@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   �\@�r����?
             .@������������������������       �                     �?�       �                   p`@@4և���?	             ,@�       �       	             �?�q�q�?             @������������������������       �                     �?�       �                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �        <            �W@�       �                    �?@��xQ�?E            �\@�       �                   �_@$�Z����?1             S@�       �                   �_@      �?             @������������������������       �                      @�       �                   q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    f@�����H�?.             R@�       �                   �m@h��@D��?-            �Q@�       �                   b@>A�F<�?             C@�       �                    @H@��a�n`�?             ?@�       �                   �k@�q�q�?             @�       �                    `@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �\@H%u��?             9@������������������������       �                      @�       �                    @J@�nkK�?             7@�       �                   P`@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@������������������������       �                     @������������������������       �                    �@@������������������������       �                     �?������������������������       �                     C@�       �       	          433�?�t����?             1@������������������������       �                     @�       �                   @i@؇���X�?	             ,@�       �                    @K@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   c@�8��8��?             (@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�                           �?Tt�ó��?#            �H@�       �                    �?      �?             C@�       �       	          ����?J�8���?             =@�       �                   `c@�q�q�?             (@������������������������       �                     @�       �                    p@����X�?             @������������������������       �                     @�       �                    �E@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    c@@�0�!��?             1@�       �                    d@      �?
             0@�       �       	          033�?��S�ۿ?	             .@������������������������       �                     (@�       �                   @`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@                        �b@���!pc�?
             &@                         �G@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @�t�b��     h�h(h+K ��h-��R�(KMKK��h_�BP       z@     P@     Pw@     @g@     `r@     @U@       @      2@       @      �?              �?       @                      1@     @r@     �P@      q@     �H@      A@      C@      9@     �A@      �?      <@      �?      0@              0@      �?                      (@      8@      @      $@      @      @      @      @       @      �?       @      �?                       @      @                      @      @              ,@              "@      @       @              �?      @               @      �?      �?              �?      �?              n@      &@      >@      "@      0@              ,@      "@      �?      @              @      �?      �?      �?                      �?      *@      @      $@      @       @       @       @                       @       @      @              �?       @       @      �?      �?      �?                      �?      �?      �?              �?      �?              @             @j@       @      @      �?      @                      �?     �i@      �?      (@      �?       @              @      �?       @               @      �?              �?       @              h@              2@      2@      @              .@      2@               @      .@      $@       @      $@      @      $@              $@      @              @              @             �S@     @Y@      &@      C@       @      @              @       @       @      @              �?       @      �?                       @      @      @@              >@      @       @      �?       @               @      �?               @              Q@     �O@      I@      :@     �@@      7@      4@      @      &@              "@      @      @      @              @      @              @              *@      4@      *@      (@      *@      "@      @      "@      @      �?              �?      @              @       @              @      @      @               @      @      @      @                      @      @                      @               @      1@      @              �?      1@       @      �?       @               @      �?              0@              2@     �B@      @      =@      @      =@      �?      �?              �?      �?               @      <@      �?      :@              0@      �?      $@              @      �?      @              @      �?      �?      �?                      �?      �?       @      �?                       @      @              &@       @       @       @       @       @              @       @       @       @                       @      @              @              F@     �s@      6@      r@      1@     @q@      @     �e@      @     �S@      @     �P@              8@      @      E@              7@      @      3@              @      @      0@       @      �?      �?              �?      �?      �?                      �?       @      .@       @      "@              @       @      @      �?              �?      @      �?                      @              @       @      *@      �?              �?      *@      �?       @              �?      �?      �?              �?      �?                      &@             �W@      &@     �Y@      &@     @P@      @      �?       @              �?      �?              �?      �?               @      P@      @      P@      @      ?@      @      8@      @       @      �?       @      �?                       @      @              @      6@       @              �?      6@      �?      @      �?                      @              .@              @             �@@      �?                      C@      @      (@      @               @      (@      �?      �?      �?                      �?      �?      &@      �?      �?      �?                      �?              $@      6@      ;@      3@      3@      $@      3@      @      @      @               @      @              @       @      �?              �?       @              @      ,@       @      ,@      �?      ,@              (@      �?       @      �?                       @      �?              �?              "@              @       @      �?       @      �?                       @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJn�GhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B(<         �                    �?�	����?R           ��@       +                   @E@J{x�%�?b           `�@                           �?�4�M�f�?B            �Y@                            P@���7�?,            �P@                          �_@0�)AU��?&            �L@������������������������       �                     C@                           �?�}�+r��?             3@       	                    �?z�G�z�?             @������������������������       �                     @
                           �J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             ,@                           �?�<ݚ�?             "@                           �?���Q��?             @������������������������       �                      @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @              	          �����X�<ݚ�?             B@                           �?r�q��?             @������������������������       �                     @������������������������       �                     �?       $                   �_@d��0u��?             >@       !       	          ����?      �?
             0@                            �?�����H�?             "@                           @K@؇���X�?             @������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @"       #                    �?և���X�?             @������������������������       �                     @������������������������       �                     @%       *                    �N@      �?             ,@&       '                    �?�z�G��?             $@������������������������       �                     @(       )                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @,       o       
             �?�������?            `|@-       ^       	          ����?����-�?`            �b@.       5                    �?�	��)��?C            �Y@/       4                    �? �Cc}�?             <@0       1       	          ����? ��WV�?             :@������������������������       �        
             .@2       3                   �Z@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �                      @6       [                   �r@���Q��?2            �R@7       D                    �?�#}7��?,            �P@8       =                   �h@��� ��?             ?@9       :                   `a@�q�q�?             "@������������������������       �                     @;       <       	          ����?      �?             @������������������������       �                     �?������������������������       �                     @>       C                   �l@���7�?             6@?       @                   �]@؇���X�?             @������������������������       �                     @A       B                    _@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     .@E       T       	          ����?)O���?             B@F       M                   0a@$��m��?             :@G       H                    �?�����H�?             2@������������������������       �                     (@I       L                    �?�q�q�?             @J       K                   g@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?N       S                    �?      �?              @O       P                    d@�q�q�?             @������������������������       �                     �?Q       R                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @U       V                    �D@z�G�z�?             $@������������������������       �                     �?W       X       	          `ff�?�����H�?             "@������������������������       �                     @Y       Z                    c@      �?              @������������������������       �                     �?������������������������       �                     �?\       ]                   �y@      �?              @������������������������       �                     @������������������������       �                     �?_       `                   �k@�r����?            �F@������������������������       �        	             1@a       j                   �o@d}h���?             <@b       c       
             �?X�<ݚ�?             "@������������������������       �                     @d       i                   Pm@�q�q�?             @e       h                   `l@z�G�z�?             @f       g                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?k       l                    @�}�+r��?             3@������������������������       �                     1@m       n       	          ���@      �?              @������������������������       �                     �?������������������������       �                     �?p       �                    @L@ȞYM�4�?�             s@q       r                   pj@���Rp�?�             m@������������������������       �        2            �S@s       �       	          pff�?�IєX�?_             c@t       }                   �b@@��9U��?S            @a@u       |                   0m@�z�N��?P            ``@v       w                    �I@t��ճC�?             F@������������������������       �                     A@x       y                    l@�z�G��?             $@������������������������       �                     @z       {                    �J@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �        7            �U@~                          �d@և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?�r����?             .@�       �                    �?���Q��?             @�       �                   `a@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                   �k@���@��?/            �R@�       �                   �`@(;L]n�?             >@�       �                    @�8��8��?	             (@������������������������       �                     &@������������������������       �                     �?������������������������       �        	             2@�       �                    c@�X���?             F@�       �                    a@��R[s�?            �A@�       �       	          @33�?��S���?             .@�       �                    �?�q�q�?             "@������������������������       �                      @�       �                    �?؇���X�?             @�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   @b@r�q��?             @������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �c@P���Q�?             4@������������������������       �                     0@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    @O@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?ȕ �&~�?�            �v@�       �                    �?x�K��?             �I@�       �                   �r@j���� �?	             1@�       �       	          ��� @r�q��?             (@������������������������       �                     $@������������������������       �                      @������������������������       �                     @�       �       	          ����?�t����?             A@�       �                   �s@D�n�3�?             3@�       �       
             �?d}h���?
             ,@�       �                   pl@8�Z$���?	             *@������������������������       �                     �?�       �                   0r@�8��8��?             (@������������������������       �                      @�       �                    b@      �?             @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    `@�r����?
             .@������������������������       �                     @�       �                    �J@�<ݚ�?             "@�       �                    �?�q�q�?             @�       �                   Pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    [@�l.�f��?�            ps@�       �                   �`@��
ц��?	             *@�       �       
             �?      �?              @������������������������       �                     @�       �                   q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�             
             �?�]z�}�?�            �r@�                          �R@��S�ۿ?�            �o@�                         (q@(�s���?�            �o@�       �                   �b@t�e�í�?�             i@�       �       	          `ff�?�*v��?~            @h@�       �                    �?4Qi0���?P            �^@�       �                   �i@h�a��?>            @X@������������������������       �        !            �G@�       �                   �Z@ףp=
�?             I@�       �                   @_@�E��ӭ�?	             2@������������������������       �                     @�       �                    Z@�q�q�?             (@�       �                    �?�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @@�       �                    �?�θ�?             :@�       �                   @e@�S����?             3@�       �                    �?�IєX�?             1@������������������������       �                     �?������������������������       �        
             0@������������������������       �                      @�       �                   �Z@և���X�?             @������������������������       �                      @�       �       	          ����?���Q��?             @������������������������       �                      @�       �                   �l@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    _@ ��PUp�?.            �Q@�       �                    �?$�q-�?
             *@�       �                    �H@�8��8��?	             (@������������������������       �                     @�       �       	          033@r�q��?             @������������������������       �                     @�       �                   �^@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �        $             M@�             	          `ff@և���X�?             @�                           �K@      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �        %            �I@            	             @�q�q�?             @������������������������       �                      @������������������������       �                     �?                         �?^����?            �E@      	                  (p@�t����?             A@������������������������       �                     6@
                        pf@�q�q�?             (@                         �?z�G�z�?             $@                        `]@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @                         I@�����H�?             "@������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KMKK��h_�B0        z@     `@     �v@     `h@      3@     �T@      @     �O@      �?      L@              C@      �?      2@      �?      @              @      �?      �?      �?                      �?              ,@       @      @       @      @               @       @      �?       @                      �?              @      0@      4@      @      �?      @                      �?      &@      3@      @      (@      �?       @      �?      @              @      �?      �?              �?      �?                       @      @      @      @                      @      @      @      @      @              @      @      @      @                      @      @             `u@      \@     �N@     �U@     �K@      H@      9@      @      9@      �?      .@              $@      �?              �?      $@                       @      >@     �F@      7@      F@      @      ;@      @      @              @      @      �?              �?      @              �?      5@      �?      @              @      �?      �?              �?      �?                      .@      3@      1@      1@      "@      0@       @      (@              @       @      @      �?              �?      @                      �?      �?      @      �?       @              �?      �?      �?      �?                      �?              @       @       @      �?              �?       @              @      �?      �?      �?                      �?      @      �?      @                      �?      @     �C@              1@      @      6@      @      @      @               @      @      �?      @      �?      �?              �?      �?                      @      �?              �?      2@              1@      �?      �?              �?      �?             �q@      9@     �k@      "@     �S@              b@      "@     ``@      @      `@      @     �D@      @      A@              @      @      @               @      @              @       @             �U@              @      @              @      @              *@       @      @       @       @       @      �?              �?       @              �?      �?      �?      �?                      �?      �?              $@              M@      0@      =@      �?      &@      �?      &@                      �?      2@              =@      .@      :@      "@      @       @      @      @               @      @      �?       @      �?       @                      �?      @              �?      @              @      �?       @              �?      �?      �?              �?      �?              3@      �?      0@              @      �?      @                      �?      @      @              @      @             �K@     0s@      4@      ?@      $@      @      $@       @      $@                       @              @      $@      8@       @      &@      @      &@       @      &@      �?              �?      &@               @      �?      @      �?      �?              �?      �?                       @      �?              @               @      *@              @       @      @       @      �?      �?      �?      �?                      �?      �?                      @     �A@     @q@      @      @      �?      @              @      �?      �?      �?                      �?      @              =@     �p@      1@     �m@      .@     �m@      .@     @g@      (@     �f@      &@      \@      @      W@             �G@      @     �F@      @      *@              @      @      @      @      @              @      @               @      �?       @                      �?              @@      @      4@      @      0@      �?      0@      �?                      0@       @              @      @               @      @       @       @              �?       @      �?                       @      �?     �Q@      �?      (@      �?      &@              @      �?      @              @      �?       @               @      �?                      �?              M@      @      @      @      �?      �?      �?      �?                      �?       @                      @             �I@       @      �?       @                      �?      (@      ?@      @      >@              6@      @       @       @       @      �?       @      �?                       @      �?               @               @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ!{�0hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK兔h~�B2         �                    �?�O(�.��?M           ��@       5                    �?��i[)f�?]           Ѐ@              
             �?4�.�A�?�            �g@                          xr@ZՏ�m|�?E            �X@                          �`@X�EQ]N�?=            �U@                          `]@�:�B��?)            �M@������������������������       �                     3@       	       	            �?      �?             D@������������������������       �                     3@
                           b@�G��l��?             5@              	          ����?j���� �?
             1@                            H@�θ�?             *@                           �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@������������������������       �                     @������������������������       �                     @������������������������       �                     ;@                          (s@      �?             (@������������������������       �                     @������������������������       �                     @                          @E@Z��:���?<            �V@                            F@�KM�]�?             3@              	          ����?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     ,@       2                    @N@r�q��?1             R@       !                    �D@��2(&�?+            �P@                            �C@և���X�?             @������������������������       �                     @������������������������       �                     @"       #                    �?�j��b�?%            �M@������������������������       �        	             (@$       '                    �?��E�B��?            �G@%       &                   pa@      �?             @������������������������       �                     @������������������������       �                     @(       )       	          ����?��p\�?            �D@������������������������       �                     <@*       /                     L@�θ�?	             *@+       .                   `@ףp=
�?             $@,       -       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @0       1                   �j@�q�q�?             @������������������������       �                     �?������������������������       �                      @3       4                   �m@      �?             @������������������������       �                     @������������������������       �                     @6       _                    �K@"YH:>�?�            �u@7       N       
             �?������?�            0p@8       =                    �?��N`.�?"            �K@9       :                   0e@�nkK�?             7@������������������������       �                     ,@;       <                   pe@�����H�?             "@������������������������       �                     �?������������������������       �                      @>       I                   0a@     ��?             @@?       @                    @B@�ՙ/�?             5@������������������������       �                     @A       H                   �q@�E��ӭ�?             2@B       C                   �[@�r����?             .@������������������������       �                     �?D       E       	          ����?@4և���?             ,@������������������������       �                     $@F       G                   0c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @J       K                   �r@"pc�
�?             &@������������������������       �                      @L       M                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @O       P                    @G@г�wY;�?            �i@������������������������       �        7            �T@Q       ^                   �g@����&!�?H            @^@R       U                   �c@0x�!���?G            �]@S       T                    �?      �?             @������������������������       �                      @������������������������       �                      @V       W                   n@�]���?E            �\@������������������������       �        $             O@X       ]                   @[@�&=�w��?!            �J@Y       Z                    �?      �?              @������������������������       �                     @[       \                    @I@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                    �F@������������������������       �                      @`       e                   �X@�L�lRT�?;            �V@a       d                    �?ףp=
�?             $@b       c                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @f       }       
             �?���Q8�?5             T@g       h                   �^@��J�fj�?            �B@������������������������       �                     @i       n       	          ����?�z�G��?             >@j       m                    �?      �?             @k       l                   0b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @o       t                    �?�θ�?             :@p       q                    �P@      �?	             0@������������������������       �                     $@r       s                    �Q@�q�q�?             @������������������������       �                      @������������������������       �                     @u       x                    �N@���Q��?             $@v       w                    �L@�q�q�?             @������������������������       �                     �?������������������������       �                      @y       z                    �P@����X�?             @������������������������       �                     @{       |       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @~       �       	          `ff�?�T|n�q�?            �E@       �                    @ףp=
�?             D@�       �                    �?�FVQ&�?            �@@������������������������       �        	             ,@�       �                   �a@�KM�]�?             3@������������������������       �                     (@�       �                   ps@����X�?             @�       �                   0b@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                   hp@����X�?             @�       �                    �?r�q��?             @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   �c@fGk�T�?�            �w@�       �                    �?�+I�9��?�            @v@�       �                    �R@ 	��p�?�             r@�       �                    �?���.�d�?�            �q@������������������������       �        $             R@�       �       	          033�?��-#���?�            �j@�       �                   �j@z�G�z�?              I@������������������������       �                    �B@�       �                     P@�θ�?
             *@�       �                   �o@�C��2(�?             &@�       �                     L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �L@H�!b	�?u            @d@�       �                   �[@DE�SA_�?F            @X@�       �                     E@      �?              @������������������������       �                     @�       �                   `_@      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                     �?�       �       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   pp@���M�??            @V@�       �                   p@ܷ��?��?)             M@�       �       	          `ff�?x�}b~|�?(            �L@�       �                    �?��hJ,�?             A@�       �                   `@      �?             @������������������������       �                     @������������������������       �                     @�       �       	          033�?@4և���?             <@�       �                   �i@���7�?             6@������������������������       �                     &@�       �                   @j@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                    b@r�q��?             @������������������������       �                     @�       �                    @H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@������������������������       �                     �?������������������������       �                     ?@������������������������       �        /            @P@�       �                   �[@�q�q�?             @������������������������       �                     @�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �`@:ɨ��?$            �P@�       �                   �\@�T|n�q�?            �E@�       �                   �Z@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �       
             �?�L���?            �B@������������������������       �                     A@������������������������       �                     @�       �                   �o@\X��t�?             7@�       �                    b@@4և���?             ,@�       �                    �H@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                   �a@�q�q�?             8@�       �       	             �?���N8�?             5@�       �                   �^@�t����?             1@������������������������       �                     @�       �                   r@"pc�
�?             &@�       �                   pd@ףp=
�?             $@�       �                    @J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �       	          033@      �?             @�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�BP       �z@     �~@     0w@     �d@     �S@     �[@      0@     �T@      $@      S@      $@     �H@              3@      $@      >@              3@      $@      &@      $@      @      $@      @      �?      @      �?                      @      "@                      @              @              ;@      @      @      @                      @      O@      =@       @      1@       @      @       @                      @              ,@      N@      (@     �L@      "@      @      @      @                      @     �J@      @      (@             �D@      @      @      @      @                      @      C@      @      <@              $@      @      "@      �?      @      �?      @                      �?      @              �?       @      �?                       @      @      @      @                      @     Pr@      L@     `m@      8@     �B@      2@      6@      �?      ,@               @      �?              �?       @              .@      1@      *@       @              @      *@      @      *@       @              �?      *@      �?      $@              @      �?              �?      @                      @       @      "@               @       @      �?              �?       @             �h@      @     �T@             �\@      @     �\@      @       @       @               @       @             @\@       @      O@             �I@       @      @       @      @              @       @               @      @             �F@                       @      M@      @@      �?      "@      �?       @      �?                       @              @     �L@      7@      5@      0@              @      5@      "@      �?      @      �?      �?              �?      �?                       @      4@      @      ,@       @      $@              @       @               @      @              @      @      �?       @      �?                       @      @       @      @              �?       @      �?                       @      B@      @      B@      @      ?@       @      ,@              1@       @      (@              @       @      @      �?              �?      @                      �?      @       @      @      �?       @      �?       @                      �?      @                      �?              @      L@     @t@      D@     �s@      4@     �p@      2@     �p@              R@      2@     @h@      $@      D@             �B@      $@      @      $@      �?       @      �?       @                      �?       @                       @       @     @c@       @     @V@       @      @              @       @       @              �?       @      �?      �?              �?      �?      �?                      �?      @     �T@      @      J@      @      J@      @      =@      @      @              @      @               @      :@      �?      5@              &@      �?      $@      �?                      $@      �?      @              @      �?      �?      �?                      �?              7@      �?                      ?@             @P@       @      @              @       @      �?              �?       @              4@      G@      @      B@      @       @               @      @              @      A@              A@      @              *@      $@      *@      �?      @      �?              �?      @              @                      "@      0@       @      0@      @      .@       @      @              "@       @      "@      �?      �?      �?      �?                      �?       @                      �?      �?      @      �?      �?      �?                      �?               @              @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KKh~�BH4         r                    �?>���i��?H           ��@       =       
             �?r|7k�?1           `@       0                   Hr@ ]�� ��?�            �v@                           �?��}� �?�            `s@              	          ����?f���M�?             ?@                           �?���Q��?
             .@������������������������       �                     @       	                    ^@      �?              @������������������������       �                     @
                           �N@���Q��?             @������������������������       �                      @������������������������       �                     @              	          pff�?      �?             0@                           �?����X�?             @                          @_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     "@       /                    �?� {��?�            pq@       "                   �a@��-��ĳ?n            �e@       !       	             �?�'F�3�?]            �b@                           �?�C��2(�?            �@@                           `@ 7���B�?             ;@                           �N@�C��2(�?             &@������������������������       �                     "@                          `^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             0@                           `^@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        H             ]@#       (                   `h@�J�4�?             9@$       '                   �g@և���X�?             @%       &                   �W@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @)       .       	          ����?�X�<ݺ?             2@*       +                    �?؇���X�?             @������������������������       �                      @,       -       	             �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �        >            @Z@1       2                   �r@R�}e�.�?              J@������������������������       �                     @3       6       
             �?�q�q�?             H@4       5                    �?և���X�?             @������������������������       �                     @������������������������       �                     @7       <                    �?��r._�?            �D@8       ;                    `@      �?             ,@9       :       	          ���@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     ;@>       Y                   �_@N� ˔x�?P            �a@?       L       	          ����?     x�?$             P@@       A                    �?�4�����?             ?@������������������������       �                     @B       I                    �?X�Cc�?             <@C       D                   Pb@��H�}�?             9@������������������������       �        	             ,@E       F                    �?"pc�
�?             &@������������������������       �                      @G       H                   �k@�q�q�?             @������������������������       �                      @������������������������       �                     �?J       K                   �r@�q�q�?             @������������������������       �                      @������������������������       �                     �?M       T       	          ����?<���D�?            �@@N       O                    �?�z�G��?             $@������������������������       �                      @P       S                    �?      �?              @Q       R                    V@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @U       V       	          ����?�nkK�?             7@������������������������       �        
             5@W       X                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?Z       c                    �?p9W��S�?,             S@[       `                    @N@Du9iH��?            �E@\       ]                     I@ ���J��?            �C@������������������������       �        
             2@^       _       	          `ffֿ���N8�?             5@������������������������       �                     �?������������������������       �                     4@a       b                   �j@      �?             @������������������������       �                      @������������������������       �                      @d       q                   �f@4���C�?            �@@e       h                    @I@l��[B��?             =@f       g                    �F@r�q��?             @������������������������       �                     �?������������������������       �                     @i       j                    �?�û��|�?             7@������������������������       �                     @k       l       	             �?�z�G��?             4@������������������������       �                     @m       p                    S@��S�ۿ?	             .@n       o                   �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                     @s       �       
             �?t�n_Y��?            z@t       �                   �b@�r�K��?j            `d@u       �                    �?�-���?F             Y@v       �                     P@և���X�?             5@w       �                    �?��.k���?             1@x       {                    @K@      �?
             0@y       z                   �a@؇���X�?             @������������������������       �                     �?������������������������       �                     @|       �                   �`@�<ݚ�?             "@}       �                    @�q�q�?             @~       �                    �?z�G�z�?             @       �                   (r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   p`@��t���?8            �S@�       �       	          `ff�?@4և���?             E@�       �                    �?ȵHPS!�?             :@������������������������       �                     �?�       �       	             �?HP�s��?             9@������������������������       �                     6@�       �                   o@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     0@�       �                   @a@V������?            �B@�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�       �                   0m@r٣����?            �@@�       �                   k@���Q��?             .@�       �                    �F@�<ݚ�?             "@������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   Pb@�q�q�?             @������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	            �?�����H�?	             2@�       �                   �a@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     ,@�       �                   Pc@p�EG/��?$            �O@������������������������       �                     &@�       �                   ``@��B����?             J@�       �                    @L@*O���?             B@�       �                    K@�c�Α�?             =@������������������������       �                      @�       �                   (p@�<ݚ�?             ;@�       �                    �C@�J�4�?             9@�       �                    @      �?             @������������������������       �                      @������������������������       �                      @�       �                   Pl@�����?             5@������������������������       �                     *@�       �       	          ����?      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?����X�?             @������������������������       �                     @�       �                   �x@      �?             @������������������������       �                      @������������������������       �                      @�       �                   pc@      �?	             0@������������������������       �                     @�       �                    �?$�q-�?             *@�       �                     @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�       �       	          ���@<��ٵ�?�            �o@�       �                   0h@`�ҕ�ļ?�            `o@�       �                   �O@��/�n�?�             o@�       �       	          ����?     ��?
             0@�       �                    �?�8��8��?             (@������������������������       �                     @�       �                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    @L@XB���?�             m@�       �                    c@�x�V�?�             g@�       �                   �b@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�o"Q9a�?            �f@�       �                   @[@�h%�M��?w            `e@�       �                    @G@؇���X�?
             ,@������������������������       �                     "@�       �                     H@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �        m            �c@������������������������       �                     $@�       �                    �L@�*/�8V�?            �G@�       �                   �`@      �?             @������������������������       �                     @������������������������       �                     @�       �                    q@������?            �D@������������������������       �                     7@�       �                    `@�����H�?
             2@������������������������       �                     �?�       �                    �?�IєX�?	             1@�       �                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     ,@�       �                    d@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@     �[@     px@      @@     �t@      2@     @r@      &@      4@      "@      @      @               @      @              @       @      @       @                      @       @      ,@       @      @       @       @       @                       @              @              "@      @      q@      @     �d@      @     @b@      @      >@      �?      :@      �?      $@              "@      �?      �?              �?      �?                      0@       @      @              @       @                      ]@      @      5@      @      @      �?      @      �?                      @       @              �?      1@      �?      @               @      �?      @              @      �?                      &@             @Z@      ,@      C@      @              $@      C@      @      @              @      @              @      A@      @      @      @       @      @                       @              @              ;@     �S@     �N@      9@     �C@      5@      $@      @              2@      $@      0@      "@      ,@               @      "@               @       @      �?       @                      �?       @      �?       @                      �?      @      =@      @      @               @      @      @      @      @              @      @                       @      �?      6@              5@      �?      �?      �?                      �?      K@      6@      D@      @      C@      �?      2@              4@      �?              �?      4@               @       @               @       @              ,@      3@      ,@      .@      @      �?              �?      @              "@      ,@      @              @      ,@      @              �?      ,@      �?      @              @      �?                      &@              @     �r@      ]@      P@     �X@      :@     �R@      (@      "@       @      "@       @       @      @      �?              �?      @               @      @       @      @      �?      @      �?       @      �?                       @               @      �?                      @              �?      @              ,@     @P@      @     �C@      @      7@      �?               @      7@              6@       @      �?       @                      �?              0@      &@      :@      @      �?      @                      �?       @      9@      @      "@       @      @      �?              �?      @              @      �?      �?              �?      �?              @       @      @              �?       @               @      �?               @      0@       @       @               @       @                      ,@      C@      9@      &@              ;@      9@      7@      *@      5@       @               @      5@      @      5@      @       @       @       @                       @      3@       @      *@              @       @      @              �?       @      �?                       @               @       @      @              @       @       @               @       @              @      (@      @              �?      (@      �?      �?      �?                      �?              &@     �m@      1@     �m@      .@     `m@      *@      &@      @      &@      �?      @              @      �?              �?      @                      @      l@       @     �f@      @      @      �?      @                      �?     `f@       @      e@       @      (@       @      "@              @       @               @      @             �c@              $@              E@      @      @      @              @      @             �C@       @      7@              0@       @              �?      0@      �?       @      �?       @                      �?      ,@              �?       @      �?                       @               @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��-]hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�9         t                   p`@TU�`��??           ��@       M                    �?B_��V��?	           P{@       2       	          ����?�L"��?�            t@       -                    �?����k��?Y            �b@              
             �?�Sb(�	�?A             [@                          �Z@z�G�z�?1             T@������������������������       �                     @                           �?؇���X�?/            @S@	       
       	            �?�<ݚ�?             "@������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     @              	          ����?�IєX�?)             Q@������������������������       �                    �A@              	          ����?<���D�?            �@@              	          hff�?      �?              @������������������������       �                     �?                           �?և���X�?             @������������������������       �                      @                           �?z�G�z�?             @                          �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     9@       &                    �?      �?             <@       !                    �L@�eP*L��?             &@                           `V@r�q��?             @                           �G@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @"       %                    \@z�G�z�?             @#       $                    d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @'       ,       	          @33�?�t����?             1@(       )                   �]@      �?             0@������������������������       �                     (@*       +                   �`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?.       1                   �X@ףp=
�?             D@/       0                    k@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @@3       J                    �Q@jه��?i            �e@4       I                    �? eD5�Ҽ?e            �d@5       8                    �?���}<S�?F            �\@6       7                    �M@�θ�?             *@������������������������       �                     $@������������������������       �                     @9       D       	          ����?�v�\�?A            �Y@:       A                    �N@���y4F�?             3@;       <                    �E@      �?             0@������������������������       �                     �?=       >                   @_@��S�ۿ?             .@������������������������       �                     &@?       @                   0j@      �?             @������������������������       �                     �?������������������������       �                     @B       C                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?E       F                    �?P��BNֱ?3            �T@������������������������       �        '            �P@G       H                   �_@     ��?             0@������������������������       �                     @������������������������       �                     *@������������������������       �                     J@K       L                   �[@�q�q�?             @������������������������       �                     @������������������������       �                      @N       g       	          033�?���N��?G             ]@O       R                    @J@�'N��?(            �N@P       Q                   �S@�C��2(�?             6@������������������������       �                      @������������������������       �                     4@S       V                    �?�n_Y�K�?            �C@T       U       
             �?8�Z$���?             *@������������������������       �                      @������������������������       �                     &@W       f       
             �?      �?             :@X       Y       
             �?�E��ӭ�?             2@������������������������       �                      @Z       e                    �?     ��?             0@[       b                    @�θ�?             *@\       ]                    �?ףp=
�?             $@������������������������       �                     �?^       a                    �L@�����H�?             "@_       `                    \@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @c       d                   c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @h       i                   @\@z�G�z�?            �K@������������������������       �        
             1@j       k                   �\@p9W��S�?             C@������������������������       �                     @l       o                   P`@4�2%ޑ�?            �A@m       n       	          ����?���Q��?             $@������������������������       �                     @������������������������       �                     @p       s                   �c@HP�s��?             9@q       r                    �? �q�q�?             8@������������������������       �                     �?������������������������       �                     7@������������������������       �                     �?u       �                    �?�P�+�?6           ~@v       �                    �?N(1����?{            @f@w       �       
             �?v ��?            �E@x       �                    �?      �?             8@y       �                    �?z�G�z�?	             .@z              	          ����?�z�G��?             $@{       ~                   �b@      �?             @|       }                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                   `T@�KM�]�?             3@������������������������       �                     �?�       �                   �b@�X�<ݺ?             2@������������������������       �        	             0@�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?��Hg���?^            �`@�       �       
             �?*-ڋ�p�?6            @S@�       �                   r@(;L]n�?             >@������������������������       �                     ;@�       �                    @F@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   ``@֭��F?�?"            �G@�       �                   �b@���Q��?             9@������������������������       �                     @�       �                    �?����X�?             5@�       �       	          ����?      �?             0@�       �                     I@���Q��?             .@�       �                   `\@���Q��?             $@�       �                   �c@      �?             @������������������������       �                     @������������������������       �                     �?�       �                     B@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �D@��2(&�?             6@������������������������       �                     �?�       �                   �i@�����?             5@�       �                   �e@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �        	             .@�       �                   `a@�8���?(             M@�       �       
             �?      �?              @������������������������       �                     @������������������������       �                      @�       �                    U@p���?!             I@�       �                    �J@�8��8��?             (@�       �       	          ����?z�G�z�?             @������������������������       �                     @�       �                   �W@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     C@�       �                    �?JD�����?�            �r@�       �                    �?��g=��?Q            @a@�       �                   @g@      �?J             `@�       �       	          ���@X�GP>��?I            �_@�       �                    �?���N8�?H            �_@�       �                    �?r�q��?
             (@�       �                   `n@�q�q�?             @�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   `l@���U�?>            �\@������������������������       �                    �J@�       �                    m@��GEI_�?"            �N@������������������������       �                      @�       �                   `p@���#�İ?!            �M@�       �       
             �?�����H�?             2@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   Hp@��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                    �D@������������������������       �                     �?������������������������       �                     �?�       �       	             �?      �?             $@������������������������       �                     @�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       
             �?���!pc�?j            �d@�       �                   Pb@      �?-            �Q@�       �       	          `ff�?�S����?             3@�       �                   �i@���!pc�?             &@������������������������       �                     @�       �                   0o@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?�"U����?!            �I@�       �                    �?��S�ۿ?	             .@������������������������       �                     ,@������������������������       �                     �?�       �                   �g@      �?             B@�       �                   �c@؇���X�?             @������������������������       �                     @�       �                   �S@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �`@�f7�z�?             =@�       �                    @@�0�!��?             1@�       �       	          ����?$�q-�?             *@������������������������       �                     �?������������������������       �                     (@�       �       	          ����?      �?             @������������������������       �                     �?�       �       	          ���@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   f@      �?             (@�       �                    d@ףp=
�?             $@������������������������       �                     @�       �                   p@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    @M@�KM�]�?=            �W@������������������������       �        /            �P@�                         �`@X�Cc�?             <@�                          @�eP*L��?             &@�                            P@      �?              @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @                        @t@������?             1@������������������������       �                     (@                         �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�t�b�])     h�h(h+K ��h-��R�(KMKK��h_�Bp       @y@     �@     �Z@     �t@     �I@     �p@     �C@     @[@     �A@     @R@      ,@     �P@      @              &@     �P@      @       @              �?      @      �?              �?      @              @      P@             �A@      @      =@      @      @      �?              @      @       @              �?      @      �?      �?      �?                      �?              @              9@      5@      @      @      @      @      �?      �?      �?              �?      �?              @              �?      @      �?      �?      �?                      �?              @      .@       @      .@      �?      (@              @      �?      @                      �?              �?      @      B@      @      @              @      @                      @@      (@      d@      $@     �c@      $@     @Z@      @      $@              $@      @              @     �W@      @      .@       @      ,@      �?              �?      ,@              &@      �?      @      �?                      @       @      �?       @                      �?      @      T@             �P@      @      *@      @                      *@              J@       @      @              @       @             �K@     �N@      F@      1@      4@       @               @      4@              8@      .@      &@       @               @      &@              *@      *@      @      *@       @              @      *@      @      $@      �?      "@              �?      �?       @      �?      @              @      �?                      @       @      �?              �?       @                      @       @              &@      F@              1@      &@      ;@      @               @      ;@      @      @      @                      @       @      7@      �?      7@      �?                      7@      �?             �r@     �f@     �J@     @_@      4@      7@      @      5@      @      (@      @      @      @      �?      �?      �?      �?                      �?       @                      @              @              "@      1@       @              �?      1@      �?      0@              �?      �?      �?                      �?     �@@     �Y@      >@     �G@      �?      =@              ;@      �?       @               @      �?              =@      2@      $@      .@      @              @      .@      @      $@      @      "@      @      @      �?      @              @      �?              @      �?              �?      @                      @              �?              @      3@      @              �?      3@       @      @       @      @                       @      .@              @     �K@       @      @              @       @              �?     �H@      �?      &@      �?      @              @      �?      �?      �?                      �?              @              C@     �n@      M@     @_@      *@      ^@       @      ^@      @      ^@      @      $@       @      @       @      �?       @               @      �?              @              @             �[@      @     �J@             �L@      @               @     �L@       @      0@       @       @      �?       @                      �?      ,@      �?      ,@                      �?     �D@                      �?              �?      @      @      @              �?      @      �?                      @      ^@     �F@     �A@     �A@      @      0@      @       @              @      @      @      @                      @               @      @@      3@      ,@      �?      ,@                      �?      2@      2@      �?      @              @      �?       @      �?                       @      1@      (@      ,@      @      (@      �?              �?      (@               @       @              �?       @      �?       @                      �?      @      "@      �?      "@              @      �?       @      �?                       @       @             @U@      $@     �P@              2@      $@      @      @      @      @      @      @      @                      @       @                      @      *@      @      (@              �?      @      �?                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�f6uhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�Bx=         �       
             �?�5�C��?P           ��@       ]                   �a@������?H           �@       *                    �?`�j���?�            �v@                           �?T��?D            �Y@                           @      �?             8@              	          ����?�z�G��?             4@������������������������       �                     @                          �`@ҳ�wY;�?	             1@	              	          ����?�8��8��?             (@
                          `[@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @       !                    @O@�:�^���?6            �S@                            �? ��WV�?&             J@                          `]@P���Q�?             D@������������������������       �                     7@                           �?�t����?             1@                          ``@@4և���?             ,@������������������������       �                     "@                           p@z�G�z�?             @������������������������       �                     @              	             �?      �?              @������������������������       �                     �?������������������������       �                     �?              	          `ff�?�q�q�?             @������������������������       �                     �?                          `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@"       #       
             �?���B���?             :@������������������������       �                     �?$       )                    �?�J�4�?             9@%       (                   �l@���|���?             &@&       '       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �        	             ,@+       4                    �?�'�=z��?�            �p@,       /                    @J@�	j*D�?             *@-       .       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?0       1                   0r@z�G�z�?	             $@������������������������       �                     @2       3                   �]@���Q��?             @������������������������       �                     @������������������������       �                      @5       \                    �R@�"�<F��?�            `o@6       W                    a@o�U��?�             o@7       F                    �?0]Z �i�?�            @m@8       ?       	          ����?�h%�M��?j            `e@9       :                   �`@`2U0*��?             9@������������������������       �        
             .@;       <                   �\@ףp=
�?             $@������������������������       �                      @=       >                    �?      �?              @������������������������       �                     �?������������������������       �                     �?@       E                    \@�1���܋?Y            @b@A       D       	             �?�8��8��?             (@B       C                    ^@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �        Q            �`@G       L                   `X@���N8�?'            �O@H       I                    @K@����X�?             @������������������������       �                     @J       K                    W@�q�q�?             @������������������������       �                     �?������������������������       �                      @M       V                    �?�h����?#             L@N       O                   �n@P�Lt�<�?             C@������������������������       �                     9@P       Q       
             �?$�q-�?             *@������������������������       �                     �?R       U                   `\@�8��8��?             (@S       T                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@������������������������       �                     2@X       [       	             �?�r����?             .@Y       Z                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@������������������������       �                      @^       s                    �?L�w�=�?[            �a@_       h                    �?�?�<��?+            @P@`       g                    �?�t����?             1@a       f       	          033@      �?             $@b       e                    �N@r�q��?             @c       d                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @i       l                   �b@      �?              H@j       k       	          hff�?r�q��?	             (@������������������������       �                      @������������������������       �                     $@m       r                    �?������?             B@n       o                     M@�IєX�?             1@������������������������       �        
             .@p       q                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     3@t       w                    @B@�EH,���?0            �R@u       v                    ]@؇���X�?             @������������������������       �                     �?������������������������       �                     @x       �                    �?�)�8��?-             Q@y       z                   Ph@      �?
             0@������������������������       �                      @{       ~                   0q@؇���X�?	             ,@|       }                    �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@       �                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          pff�?��B����?#             J@������������������������       �                     @�       �                   g@(옄��?             G@�       �                     P@X��ʑ��?            �E@�       �       	             �?�G�z��?             D@�       �                   �i@      �?
             0@������������������������       �                     �?�       �                    �?z�G�z�?	             .@�       �                   b@r�q��?             (@������������������������       �                     @�       �                   @b@����X�?             @������������������������       �                     �?�       �                    c@r�q��?             @�       �                    _@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          @33�?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   �l@�q�q�?             8@�       �                   f@�z�G��?             $@�       �                   �c@      �?             @������������������������       �                      @�       �       	          `ff@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       
             �?d}h���?	             ,@������������������������       �                     @������������������������       �                     &@������������������������       �                     @������������������������       �                     @�       �                    P@�}�	���?           �y@�       �                    Z@������?!            �I@�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �?:	��ʵ�?            �F@�       �                    @M@�ՙ/�?             5@�       �                    �J@ףp=
�?             $@������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?���|���?	             &@�       �                    �?      �?             @�       �       	             п      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   `V@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     8@�                          �?ıD���?�            �v@�             	          033@�2bC�?�            t@�       �                    �?��6r1-�?�            �s@�       �                    �?r�q��?2            �V@�       �                   �a@�q�q�?             8@������������������������       �                     (@�       �                   f@�q�q�?	             (@�       �                    �H@z�G�z�?             $@������������������������       �                     @�       �       	          @33�?�q�q�?             @�       �                   �`@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   pc@��IF�E�?%            �P@�       �       	          hff�?@��8��?             H@������������������������       �                    �G@������������������������       �                     �?�       �                   �c@�q�q�?             2@������������������������       �                     @�       �                    ]@z�G�z�?
             .@������������������������       �                     �?�       �                   �b@؇���X�?	             ,@�       �                   �_@$�q-�?             *@�       �                    _@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                     �?�       �                    �?���U�?�            �l@�       �                    @�KM�]�?             C@�       �                   �`@�FVQ&�?            �@@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�g�y��?             ?@�       �                   �a@��S�ۿ?	             .@������������������������       �                     *@�       �                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             0@�       �                   �a@���Q��?             @������������������������       �                      @������������������������       �                     @�                           @ r���?�            �g@�       �                    �?0m��5!�?{            �f@�       �       	            �?�{���l�?h            �c@�       �                    �O@`��(�?Y            �`@�       �                    �?@M^l���?W            �`@�       �                   @[@ �|ك�?P            �^@�       �                    �?@4և���?             ,@������������������������       �                      @�       �                   @Z@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        H            @[@������������������������       �                     $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�C��2(�?             6@�       �                    �?r�q��?	             (@������������������������       �                     @�       �                   �_@���Q��?             @�       �                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     8@������������������������       �                     "@������������������������       �                     @                         �?�Q����?             D@                        (p@d��0u��?             >@                         �L@�<ݚ�?             2@            	             �?���|���?             &@                         b@      �?              @������������������������       �                     @	      
                   @K@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         �?�q�q�?             (@������������������������       �                      @            	          ����?      �?             $@                        �r@����X�?             @                         �?r�q��?             @                        `e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KMKK��h_�B�       �y@     �@      U@     `z@      C@     �t@      9@     @S@      2@      @      ,@      @      @              &@      @      &@      �?      @      �?              �?      @               @                      @      @              @     �Q@       @      I@       @      C@              7@       @      .@      �?      *@              "@      �?      @              @      �?      �?              �?      �?              �?       @              �?      �?      �?      �?                      �?              (@      @      5@      �?              @      5@      @      @      @       @               @      @                      @              ,@      *@     `o@      @      "@       @      �?       @                      �?       @       @              @       @      @              @       @              "@     @n@      @     @n@      @     �l@       @      e@      �?      8@              .@      �?      "@               @      �?      �?      �?                      �?      �?      b@      �?      &@      �?      @              @      �?                      @             �`@      @      N@       @      @              @       @      �?              �?       @              �?     �K@      �?     �B@              9@      �?      (@              �?      �?      &@      �?       @      �?                       @              "@              2@       @      *@       @      @              @       @                      $@       @              G@     �W@       @     �L@      @      (@      @      @      @      �?       @      �?       @                      �?      @                      @              @      @     �F@       @      $@       @                      $@      �?     �A@      �?      0@              .@      �?      �?      �?                      �?              3@      C@     �B@      �?      @      �?                      @     �B@      ?@      (@      @               @      (@       @      &@      �?              �?      &@              �?      �?              �?      �?              9@      ;@              @      9@      5@      6@      5@      6@      2@      (@      @              �?      (@      @      $@       @      @              @       @              �?      @      �?       @      �?       @                      �?      @               @      �?              �?       @              $@      ,@      @      @      �?      @               @      �?      �?              �?      �?              @              @      &@      @                      &@              @      @             �t@      U@      (@     �C@      @       @      @                       @       @     �B@       @      *@      �?      "@              @      �?      @              @      �?              @      @      �?      @      �?      �?      �?                      �?               @      @      �?              �?      @                      8@     �s@     �F@     pr@      :@     pr@      7@     �R@      .@      0@       @      (@              @       @       @       @              @       @      @       @      @              @       @                      �?       @             �M@      @     �G@      �?     �G@                      �?      (@      @              @      (@      @              �?      (@       @      (@      �?      @      �?      @                      �?      "@                      �?     �k@       @      A@      @      ?@       @      �?      �?      �?                      �?      >@      �?      ,@      �?      *@              �?      �?              �?      �?              0@              @       @               @      @             @g@      @      f@      @      c@      @     �`@       @     �`@      �?     �^@      �?      *@      �?       @              @      �?      @                      �?     @[@              $@              �?      �?      �?                      �?      4@       @      $@       @      @              @       @      �?       @               @      �?               @              $@              8@              "@                      @      5@      3@      &@      3@      @      ,@      @      @      @      @      @              �?      @              @      �?                      @              @      @      @       @              @      @      @       @      @      �?      �?      �?              �?      �?              @                      �?              @      $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B88         �                    �?��/.��?A           ��@       M       	          033�?�B��T�?8           �}@       $       
             �?h��7���?�            `i@                          0l@\�t��Y�?B            �Y@                          �h@0�z��?�?*             O@������������������������       �        !             I@                          �_@�8��8��?	             (@������������������������       �                      @	       
                   `^@      �?             @������������������������       �                      @                           �J@      �?              @������������������������       �                     �?������������������������       �                     �?                           �?���� �?            �D@                          `a@��
ц��?             *@              	          ����?r�q��?             @                           c@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                            M@����X�?             @              	            �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @                           �?؇���X�?             <@                          �c@      �?	             0@              	          ����?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                      @        #                    b@      �?             (@!       "       	          833�?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @%       <                   �b@�JY�8��?A             Y@&       +                    �?      �?(             N@'       (                    �L@և���X�?             @������������������������       �                      @)       *                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?,       -                    U@ {��e�?#            �J@������������������������       �                     @.       3                    �?�J�4�?!             I@/       2                    �E@���H��?             E@0       1                   @_@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     A@4       5                   �Z@      �?              @������������������������       �                     �?6       ;                   �Z@����X�?             @7       :       	             �?      �?             @8       9                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @=       J                   ``@�G�z��?             D@>       I                   `u@�	j*D�?             :@?       @                   �g@ �o_��?             9@������������������������       �                     @A       D                    �I@�q�q�?             5@B       C                   pc@      �?              @������������������������       �                      @������������������������       �                     @E       H                    �?$�q-�?             *@F       G                   d@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?K       L                    b@����X�?             ,@������������������������       �                     $@������������������������       �                     @N       i                    �?���P��?�            0q@O       h                    �Q@��a�n`�?)             O@P       W       	          ����?F�4�Dj�?(            �M@Q       V                   pr@      �?             0@R       S       
             �?�C��2(�?             &@������������������������       �                     @T       U                   �`@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @X       a                    �?X�EQ]N�?            �E@Y       Z                   Pj@      �?              @������������������������       �                     �?[       \                    �?����X�?             @������������������������       �                      @]       `                    �?���Q��?             @^       _                   �u@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?b       g                    �? >�֕�?            �A@c       d                    ]@�r����?	             .@������������������������       �                     "@e       f                   �Z@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     4@������������������������       �                     @j       s                    @G@����Q8�?�            �j@k       p                    �?r�q��?             8@l       o                   �e@�����?             5@m       n                    e@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �        
             (@q       r                    ^@�q�q�?             @������������������������       �                      @������������������������       �                     �?t       �                    �?�J�-/��?z            �g@u       �                   �a@ȵHPS!�?             :@v       {                   �q@     ��?	             0@w       z                   h@$�q-�?             *@x       y                   @_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@|       }                    �?�q�q�?             @������������������������       �                     �?~                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �       
             �?0�`G�r�?k            `d@�       �       	          033@`����֜?]            �a@������������������������       �        F            �Y@�       �                   �_@@-�_ .�?            �B@�       �                   �p@      �?              @�       �       	          `ff
@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     =@�       �                   �`@�LQ�1	�?             7@������������������������       �        	             .@�       �                   `W@      �?              @������������������������       �                     @������������������������       �                     @�       �                    �K@x��}�?	           �{@�       �                    @G@�q��/��?�            @q@�       �                   �c@PF��t<�?N            �_@�       �                   �`@�θ�?             *@������������������������       �                      @�       �                    @�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�       �       	          033@�Ru߬Α?H            �\@������������������������       �        G            @\@������������������������       �                     �?�       �                   `c@��H�&p�?]            �b@�       �                   �`@�r����?
             .@������������������������       �                     (@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �`@p^H�&m�?S            �`@�       �                    �H@hl �&�?:             W@�       �                    �?�C��2(�?             6@������������������������       �                     &@�       �       
             �?"pc�
�?             &@�       �                    �?�q�q�?             @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    `@`����֜?+            �Q@������������������������       �                      J@�       �                    ^@�X�<ݺ?             2@������������������������       �                     �?������������������������       �        
             1@�       �       
             �?���N8�?             E@�       �                   �d@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�       �                   �f@      �?             @@������������������������       �                     ?@������������������������       �                     �?�       �                    �?z�^��?^            �d@�       �       
             �?r�0?��?@            �Z@�       �                    �?f�<�>��?$            �M@�       �                   �c@�xGZ���?            �A@�       �       	          033�?П[;U��?             =@�       �                   �a@r�q��?             8@�       �                    @ҳ�wY;�?             1@�       �                   �`@��
ц��?             *@�       �                    Y@�eP*L��?
             &@������������������������       �                      @�       �                    �?�q�q�?	             "@������������������������       �                     @�       �                    �?���Q��?             @�       �                    �?      �?             @�       �                   @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @����X�?             @�       �                    �N@      �?             @������������������������       �                     �?�       �                   �b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   0a@�q�q�?             8@�       �                   �s@�KM�]�?             3@������������������������       �        	             .@�       �                   `c@      �?             @������������������������       �                      @������������������������       �                      @�       �                   �o@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   ``@�8��8��?             H@������������������������       �                     7@�       �                    �?�J�4�?             9@������������������������       �                     (@�       �                   �`@�	j*D�?
             *@������������������������       �                      @�       �       	          ����?"pc�
�?             &@�       �                   `c@���Q��?             @�       �                     M@      �?             @������������������������       �                     �?�       �                   @c@�q�q�?             @������������������������       �                     �?�       �                    d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �b@�^���U�?            �L@�       �                   �\@�θ�?            �C@�       �                   �Z@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �`@��hJ,�?             A@������������������������       �                     2@�       �                   �`@     ��?             0@������������������������       �                     &@������������������������       �                     @�                          `a@�E��ӭ�?
             2@�       �       	          `ff@      �?             $@�       �                   �`@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KMKK��h_�B       P{@     ~@     @Y@     �w@     �R@      `@      (@     �V@      �?     �N@              I@      �?      &@               @      �?      @               @      �?      �?              �?      �?              &@      >@      @      @      @      �?      �?      �?      �?                      �?      @               @      @       @      @              @       @                       @      @      8@      �?      .@      �?      @              @      �?                       @      @      "@      @      @              @      @                      @     �O@     �B@     �F@      .@      @      @       @              �?      @              @      �?              E@      &@              @      E@       @     �B@      @      @      @              @      @              A@              @      @              �?      @       @       @       @       @      �?       @                      �?              �?      @              2@      6@       @      2@      @      2@              @      @      ,@      @       @               @      @              �?      (@      �?      @      �?                      @              @      �?              $@      @      $@                      @      :@      o@      ,@      H@      &@      H@      @      $@      �?      $@              @      �?      @              @      �?              @              @      C@      @      @      �?               @      @               @       @      @       @       @       @                       @              �?       @     �@@       @      *@              "@       @      @       @                      @              4@      @              (@      i@      @      4@       @      3@       @      @              @       @                      (@       @      �?       @                      �?       @     �f@      @      7@      @      *@      �?      (@      �?      @              @      �?                      "@       @      �?      �?              �?      �?      �?                      �?              $@      @     �c@       @     @a@             �Y@       @     �A@       @      @       @      �?       @                      �?              @              =@      @      4@              .@      @      @      @                      @      u@      Z@     �n@      >@     �^@      @      $@      @               @      $@      �?      $@                      �?     @\@      �?     @\@                      �?     �^@      :@       @      *@              (@       @      �?       @                      �?     @^@      *@     @V@      @      4@       @      &@              "@       @      �?       @      �?      �?              �?      �?                      �?       @             @Q@      �?      J@              1@      �?              �?      1@              @@      $@      �?      "@              "@      �?              ?@      �?      ?@                      �?     �V@     �R@      Q@     �C@      8@     �A@      3@      0@      *@      0@      *@      &@      &@      @      @      @      @      @       @              @      @              @      @       @      @      �?      �?      �?              �?      �?               @                      �?       @              @               @      @       @       @              �?       @      �?              �?       @                      @              @      @              @      3@       @      1@              .@       @       @       @                       @      @       @      @                       @      F@      @      7@              5@      @      (@              "@      @               @      "@       @      @       @       @       @              �?       @      �?      �?              �?      �?              �?      �?              �?              @              6@     �A@      "@      >@      @      �?              �?      @              @      =@              2@      @      &@              &@      @              *@      @      @      @      @      @      @                      @               @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJdb.hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B�4         p       	          ����?x��X���?N           ��@       A                    �?}���?2            ~@                          �a@      �?~             h@              
             �?�j��b�?!            �M@������������������������       �                     D@              	          ����?�����?             3@       
                   �]@      �?             (@       	                   e@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @       ,                    �J@��rq���?]            �`@       !                    �?4�B��?5            �R@              
             �?x��}�?)            �K@                           @J@�θ�?             *@                           Z@�C��2(�?
             &@������������������������       �                     �?������������������������       �        	             $@������������������������       �                      @                           �?@4և���?             E@                          �i@      �?              @������������������������       �                     �?                           @F@؇���X�?             @������������������������       �                     �?������������������������       �                     @                            @D@г�wY;�?             A@                          �e@r�q��?             @������������������������       �                     @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     <@"       '                    �H@D�n�3�?             3@#       $                   �`@      �?             (@������������������������       �                      @%       &                   �a@      �?             @������������������������       �                     @������������������������       �                     �?(       )                   n@����X�?             @������������������������       �                     @*       +                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @-       <                    �?6�iL�?(            �M@.       /                   �h@�P�*�?             ?@������������������������       �                     @0       1                    @M@�	j*D�?             :@������������������������       �                      @2       ;                    �?X�<ݚ�?             2@3       6                    �?�q�q�?             (@4       5                    �N@���Q��?             @������������������������       �                     @������������������������       �                      @7       :       	          ����?؇���X�?             @8       9                    @O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @=       >       
             �? �Cc}�?             <@������������������������       �                     5@?       @                    �?և���X�?             @������������������������       �                     @������������������������       �                     @B       E                    I@<�&9�?�             r@C       D       
             �?p�ݯ��?             3@������������������������       �                     (@������������������������       �                     @F       _                   �a@H�S[��?�            �p@G       Z       
             �?h�lI	��?�            �k@H       S                    �K@��J�fj�?            �B@I       R                    �?8^s]e�?             =@J       K                    �?�θ�?             :@������������������������       �                     *@L       M                    �?��
ц��?             *@������������������������       �                     @N       Q                    �?�q�q�?             "@O       P                     C@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @T       U       	          ����?      �?              @������������������������       �                     @V       Y                    �?      �?             @W       X                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @[       \                    �O@0�z��?�?s            @g@������������������������       �        m             f@]       ^                   Pc@�z�G��?             $@������������������������       �                     @������������������������       �                     @`       a                    �?     ��?             H@������������������������       �                     *@b       o                    �?և���X�?            �A@c       d                    @J@      �?             @@������������������������       �        
             (@e       n                   �p@���Q��?
             4@f       i                    �?�n_Y�K�?             *@g       h                    �O@���Q��?             @������������������������       �                     @������������������������       �                      @j       k                    �?      �?              @������������������������       �                     @l       m                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @q       �                    �?`A6�S�?           @{@r       �                    �?�eP*L��?0            @S@s       �                   �e@�X����?             F@t                           �?      �?             D@u       z       	             �?     ��?             0@v       w                    �O@؇���X�?             @������������������������       �                     @x       y                    �?      �?              @������������������������       �                     �?������������������������       �                     �?{       ~       	          `ff@�����H�?             "@|       }                   �`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   `^@      �?             8@�       �                   `c@և���X�?             @�       �                   @_@���Q��?             @�       �                    @H@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �        
             1@������������������������       �                     @�       �                   `X@6YE�t�?            �@@������������������������       �                      @�       �       
             �?��a�n`�?             ?@�       �                   �p@z�G�z�?	             .@������������������������       �                     &@�       �                     @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@�       �                    f@�["���?�            pv@�       �                   �b@�G�V�e�?�            @u@�       �                    �?��OoN��?�            �r@�       �                   �U@�8���?�             m@������������������������       �                     �?�       �       
             �?���N8�?�            �l@�       �                    �R@P�	Q��?�            �h@�       �                   �z@ ���4�?�            �h@�       �       	          ����? ����?�            `h@�       �                   �[@`�(c�?>            �X@�       �                    �?z�G�z�?
             .@�       �                   �^@և���X�?             @������������������������       �                      @�       �       	             �?���Q��?             @�       �                    b@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �        4            �T@������������������������       �        B            @X@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                   Pv@     ��?             @@�       �       	          033�?��� ��?             ?@������������������������       �                     7@�       �                   �b@      �?              @�       �                   @`@�q�q�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �       	           33@��&����?/            @P@�       �       
             �?���N8�?.            �O@�       �                    �?�iʫ{�?&            �J@�       �       	          `ff�?���!pc�?             6@�       �       	          ����?��
ц��?             *@�       �                    �?�<ݚ�?             "@�       �                    @I@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                    Y@��a�n`�?             ?@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   P`@h�����?             <@�       �                   �_@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     1@�       �                    d@���Q��?             $@������������������������       �                     @�       �                   �_@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �d@�lg����?            �E@�       �                    �?���Q��?             9@�       �                   �c@�z�G��?             $@�       �                   �Y@؇���X�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �M@z�G�z�?             .@������������������������       �                     �?�       �                    �L@؇���X�?
             ,@������������������������       �                     @�       �       
             �?����X�?             @������������������������       �                      @������������������������       �                     @�       �                    @F@�X�<ݺ?
             2@�       �                   �e@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@�       �                    �?�S����?	             3@�       �                    @�����H�?             2@������������������������       �                     @�       �                   �m@"pc�
�?             &@�       �       	          ���@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KK�KK��h_�B       0z@     0@     �s@     �d@      R@      ^@      @     �J@              D@      @      *@      @      @      @      �?      @                      �?              @              @     �P@     �P@      I@      8@      E@      *@      @      $@      �?      $@      �?                      $@       @             �C@      @      @       @              �?      @      �?              �?      @             �@@      �?      @      �?      @              �?      �?              �?      �?              <@               @      &@      @      "@               @      @      �?      @                      �?      @       @      @              �?       @      �?                       @      0@     �E@      *@      2@      @               @      2@               @       @      $@       @      @       @      @              @       @              @      �?       @      �?       @                      �?      @                      @      @      9@              5@      @      @              @      @             �n@      G@      @      (@              (@      @             �m@      A@     �i@      3@      5@      0@      4@      "@      4@      @      *@              @      @      @              @      @      @       @               @      @                      @              @      �?      @              @      �?      @      �?      �?      �?                      �?               @     �f@      @      f@              @      @      @                      @     �@@      .@      *@              4@      .@      4@      (@      (@               @      (@       @      @       @      @              @       @              @       @      @              �?       @               @      �?                      @              @     �Y@     �t@      E@     �A@      ,@      >@      $@      >@      @      "@      @      �?      @              �?      �?      �?                      �?      �?       @      �?      @      �?                      @              @      @      5@      @      @      @       @       @       @               @       @              �?                       @              1@      @              <@      @               @      <@      @      (@      @      &@              �?      @              @      �?              0@             �N@     �r@     �F@     pr@      =@     �p@      (@     �k@      �?              &@     �k@      @      h@      @      h@      @      h@      @     �W@      @      (@      @      @               @      @       @      �?       @      �?                       @       @                       @             �T@             @X@       @      �?       @                      �?      �?              @      ;@      @      ;@              7@      @      @       @      @       @      �?              �?       @                      @       @              �?              1@      H@      .@      H@      "@      F@      @      0@      @      @       @      @       @      �?       @                      �?              @      @                      "@      @      <@       @      �?       @                      �?      �?      ;@      �?      $@              $@      �?                      1@      @      @              @      @      �?              �?      @               @              0@      ;@      .@      $@      @      @      �?      @      �?      �?      �?                      �?              @       @      �?       @                      �?      (@      @              �?      (@       @      @              @       @               @      @              �?      1@      �?      @      �?                      @              ,@      0@      @      0@       @      @              "@       @      @       @      @                       @      @                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJn
4hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B9         �                    �?��e�B��?<           ��@       -       	          ����?���F@�?#           �}@                          �_@�������?d            `c@              	          ����?`���i��?             F@                           �?������?             B@������������������������       �                     <@              	             �      �?              @������������������������       �                     �?	                           �F@؇���X�?             @
                          �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @              
             �?P7Z�U��?G            �[@              	          ����?d,���O�?!            �I@������������������������       �                    �A@                           �?     ��?
             0@                           �?؇���X�?             @������������������������       �                     @������������������������       �                     �?                          �p@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @       $                    �?��0u���?&             N@                          �_@p�ݯ��?             3@                           @I@      �?              @������������������������       �                     @                           �?      �?             @������������������������       �                     �?������������������������       �                     @        #                    �?�eP*L��?             &@!       "                    �M@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @%       &                   �k@,���i�?            �D@������������������������       �                     3@'       (                   pc@�GN�z�?             6@������������������������       �        
             0@)       ,       	          ����?r�q��?             @*       +                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?.       K                    �?��T\��?�            �s@/       J                   pe@ٜSu��?*            @Q@0       ?                   �`@.��<�?(            �P@1       2                    @H@4���C�?            �@@������������������������       �                     "@3       >       
             �?�q�q�?             8@4       7                    �?���|���?             6@5       6                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?8       9                   �[@��S���?	             .@������������������������       �                     @:       =                    @P@�q�q�?             (@;       <       	             �?�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @@       I                    �?l��\��?             A@A       F                    �?z�G�z�?
             .@B       E       	          033@�����H�?             "@C       D                    b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @G       H       
             �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     3@������������������������       �                      @L       Q                    Z@j��pX�?�             o@M       N                   Pd@X�<ݚ�?             "@������������������������       �                     @O       P                   �b@z�G�z�?             @������������������������       �                     @������������������������       �                     �?R       q                   �b@X�aC�U�?�            �m@S       X                   �X@ d���W�?j            @f@T       W       	             �?"pc�
�?             &@U       V                   @^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @Y       h                    _@��Q���?d            �d@Z       [                    �F@�C��2(�?             F@������������������������       �        	             0@\       g                   pp@؇���X�?             <@]       b                   �`@z�G�z�?             4@^       _                   �^@      �?             0@������������������������       �                     &@`       a                     L@���Q��?             @������������������������       �                      @������������������������       �                     @c       d                   a@      �?             @������������������������       �                     �?e       f       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @i       j       	          033�? �|ك�?H            �^@������������������������       �        '             Q@k       l                    @M@ �Jj�G�?!            �K@������������������������       �                     =@m       p                    �M@ ��WV�?             :@n       o                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     7@r       �       	          ����?\#r��?'            �N@s       ~       
             �?�<ݚ�?             ;@t       w                     F@r�q��?             8@u       v                    �?      �?             @������������������������       �                      @������������������������       �                      @x       }                    u@ףp=
�?             4@y       |                    �H@�}�+r��?             3@z       {       	             �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             .@������������������������       �                     �?       �                   �c@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     A@�       �                    @K@$09����?           �{@�       �       	          ����?\5��P�?�            pq@�       �                    �?8�W���?�            `j@�       �                    �?���ؑ�?}            �h@�       �                    @�?�|�?v             g@�       �                   �~@�x�E~�?q            @f@�       �                    @H@P����?p             f@������������������������       �        G            �Z@�       �                    f@hA� �?)            �Q@�       �                   `]@��.N"Ҭ?(            @Q@�       �       
             �?ףp=
�?	             4@������������������������       �                      @������������������������       �                     2@������������������������       �                    �H@������������������������       �                     �?������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     @�       �                   �h@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?      �?             (@������������������������       �                     �?�       �                   �^@"pc�
�?             &@�       �                   �[@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	          @33�?X�Cc�?             ,@�       �       
             �?�q�q�?	             (@������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                    �?�v:���?)             Q@�       �       	          ����?      �?
             0@�       �                   `b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     &@�       �                   �[@��WV��?             J@�       �                    �?      �?              @�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �F@�zv�X�?             F@�       �                   @_@���N8�?             5@�       �                    @�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     $@�       �                    �?8����?             7@�       �                   �]@��S���?             .@������������������������       �                     @�       �       	          ����?�q�q�?
             (@������������������������       �                     @�       �                   �_@����X�?             @�       �                    @�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?É`���?h            �d@�       �                    �?ҳ�wY;�?N            �]@�       �                   �b@��S���?             >@�       �                   `_@������?             .@�       �                   `]@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       	          ����?ףp=
�?             $@������������������������       �                     @�       �                   �k@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?z�G�z�?	             .@�       �                    �N@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?\{��)x�?:            @V@�       �                   �p@     ��?)             P@�       �       	            �?�%^�?            �E@�       �       
             �?�n`���?             ?@������������������������       �                     @�       �                   �b@ ��WV�?             :@������������������������       �                     9@������������������������       �                     �?�       �                   o@�q�q�?	             (@�       �                    @�<ݚ�?             "@������������������������       �                     @�       �                    �O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �t@���N8�?             5@������������������������       �        	             1@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       
             �?� �	��?             9@�       �                    @O@d}h���?             ,@�       �                    @L@�����H�?             "@�       �                    _@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    `P@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       	          (33�?���!pc�?             &@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   `k@      �?             H@������������������������       �        
             5@�       �                   l@�����H�?             ;@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?�             
             �?HP�s��?             9@             	          ����? �q�q�?             8@                        `n@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     .@������������������������       �                     �?�t�b�w     h�h(h+K ��h-��R�(KMKK��h_�BP       �y@     �@     @W@     �w@     �L@     �X@      �?     �E@      �?     �A@              <@      �?      @              �?      �?      @      �?      �?              �?      �?                      @               @      L@     �K@      *@      C@             �A@      *@      @      @      �?      @                      �?      @       @      @                       @     �E@      1@      @      (@      �?      @              @      �?      @      �?                      @      @      @      @      @      @                      @       @              B@      @      3@              1@      @      0@              �?      @      �?      @      �?                      @              �?      B@     �q@      3@      I@      1@      I@      ,@      3@              "@      ,@      $@      ,@       @      @      �?      @                      �?       @      @              @       @      @       @      �?       @                      �?              @               @      @      ?@      @      (@      �?       @      �?      �?      �?                      �?              @       @      @              @       @                      3@       @              1@     �l@      @      @              @      @      �?      @                      �?      *@     @l@      @     `e@       @      "@       @      �?              �?       @                       @      @     @d@      @      D@              0@      @      8@      @      0@       @      ,@              &@       @      @       @                      @       @       @      �?              �?       @      �?                       @               @      �?     �^@              Q@      �?      K@              =@      �?      9@      �?       @               @      �?                      7@      @     �K@      @      5@      @      4@       @       @       @                       @       @      2@      �?      2@      �?      @      �?                      @              .@      �?               @      �?       @                      �?              A@     t@     @_@      n@      C@     �h@      *@     �g@       @     �f@      @     �e@      @     �e@      @     �Z@             �P@      @     �P@       @      2@       @               @      2@             �H@                      �?              �?      @      �?      @               @      �?              �?       @              "@      @              �?      "@       @      @       @      @                       @      @              "@      @      @      @              @      @               @             �E@      9@      ,@       @      @       @      @                       @      &@              =@      7@       @      @       @      @              @       @                      @      ;@      1@      4@      �?      $@      �?      $@                      �?      $@              @      0@      @       @              @      @      @      @               @      @       @      �?      �?      �?              �?      �?              �?                      @               @      T@     �U@     @S@      E@      ,@      0@      &@      @       @      @       @                      @      "@      �?      @              @      �?              �?      @              @      (@       @      &@              &@       @              �?      �?              �?      �?             �O@      :@      J@      (@      @@      &@      9@      @              @      9@      �?      9@                      �?      @      @      @       @      @              �?       @               @      �?                      @      4@      �?      1@              @      �?      @                      �?      &@      ,@      @      &@      �?       @      �?       @      �?                       @              @       @      @       @                      @       @      @      @               @      @       @                      @      @     �F@              5@      @      8@      �?      �?      �?                      �?       @      7@      �?      7@      �?       @      �?                       @              .@      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJU�\hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B(5         �                    �L@�LT ���?8           ��@       M       
             �?R��@�?h           ��@       F                   �a@x��6Y�?�            �p@       +                    �?�+e�X�?�             i@                           �?@v�禺�?T            �`@                          �Z@���|���?             6@������������������������       �                     �?                          @a@�q�q�?             5@	                           �?�����H�?             "@
                            J@؇���X�?             @                           �H@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @                           �?      �?             (@                           ^@      �?             @������������������������       �                     @������������������������       �                     @                           a@      �?             @              	          033�?      �?             @                           �I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @       &                    @L@���7�?G            �[@                          �^@p� V�?B            �Y@������������������������       �        #            �K@       %                   �\@ �q�q�?             H@                            _@r�q��?             (@������������������������       �                     �?!       $       	             �?�C��2(�?
             &@"       #       	             �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     B@'       (                    e@և���X�?             @������������������������       �                      @)       *                   �_@���Q��?             @������������������������       �                      @������������������������       �                     @,       3                    a@�������?,             Q@-       0                   �X@�S����?             3@.       /                    �?���Q��?             @������������������������       �                     @������������������������       �                      @1       2       
             �?@4և���?
             ,@������������������������       �                     �?������������������������       �        	             *@4       E                    �?���Q �?             �H@5       >                   0e@���X�K�?            �F@6       7                    T@�r����?             >@������������������������       �                      @8       =                    @L@@4և���?             <@9       :                   0a@ 7���B�?             ;@������������������������       �                     7@;       <                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �??       D                    �?���Q��?             .@@       A                    �?�eP*L��?             &@������������������������       �                     @B       C                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @G       L                    �?     ��?&             P@H       I                   Pt@�����H�?             "@������������������������       �                     @J       K                    @H@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        !            �K@N       Y                   @E@�	L �F�?�            `s@O       X                   `a@���y4F�?             3@P       S                    \@X�<ݚ�?             "@Q       R                    @B@      �?             @������������������������       �                     �?������������������������       �                     @T       W       	             �?z�G�z�?             @U       V                   `^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@Z       m                   �]@,���$�?�            0r@[       l                    ]@��[�8��?            �I@\       c                    �?��0{9�?            �G@]       ^                   c@��
ц��?             *@������������������������       �                     @_       b                    �G@؇���X�?             @`       a                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @d       k                   @[@г�wY;�?             A@e       f                    @G@      �?             0@������������������������       �                      @g       j                    c@      �?              @h       i                   �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     2@������������������������       �                     @n       y                    �? �q�q�?�             n@o       t                    �?���5��?#            �L@p       q                   �n@����?�?            �F@������������������������       �                     =@r       s                   po@      �?             0@������������������������       �                     �?������������������������       �                     .@u       x       	             �?      �?             (@v       w                    `@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @z       �       	            �?��v$���?s            �f@{       |                    �?@=��?`            �c@������������������������       �                    �E@}       �                    �?@���a��?C            �\@~       �       	          ����? ��PUp�?*            �Q@       �                    @L@@	tbA@�?(            @Q@������������������������       �        &             P@�       �                    c@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     F@�       �                    _@HP�s��?             9@�       �       	          ����?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     2@�       �                    �?������?�            �u@�       �       
             �?����*��?!            �M@�       �                    b@r�q��?             >@�       �                    �?X�Cc�?             ,@������������������������       �                      @�       �                    @P@r�q��?             @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@�       �                    �?>���Rp�?             =@�       �                   p@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     5@�       �       
             �?H~��D
�?�            �q@�       �                    �?=�Ѝ;�?}            �i@�       �                    �?,N�_� �?X            �b@������������������������       �                     B@�       �       
             �?4և����?@             \@�       �                   �^@�t����?
             1@�       �                    �?����X�?             @������������������������       �                      @�       �                   `c@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     $@�       �       	          033�?�}�+r��?6            �W@�       �                   �`@,���i�?            �D@�       �                   �_@     ��?             0@������������������������       �                     "@�       �                    `@����X�?             @������������������������       �                      @�       �       	             �?���Q��?             @������������������������       �                     �?�       �                   �`@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     9@������������������������       �                     K@�       �                   �a@�c�Α�?%             M@�       �                   �a@$G$n��?            �B@�       �                    �?���7�?             6@�       �                   `[@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     .@�       �                   �[@������?	             .@������������������������       �                     @������������������������       �                     &@�       �                    `P@�G��l��?             5@�       �       	          ����?�	j*D�?             *@������������������������       �                     @������������������������       �                     "@�       �                   �Z@      �?              @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   �]@V�K/��?2            �S@�       �                   �\@�8��8��?             (@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@�       �                   `Q@���`��?+            �P@�       �                    �?���N8�?             5@�       �                   @e@      �?             $@�       �                    �?      �?              @������������������������       �                     @�       �                   �V@���Q��?             @������������������������       �                      @�       �                   �]@�q�q�?             @������������������������       �                     �?�       �                   `_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                    �?�I� �?             G@�       �                    @     ��?             @@�       �                   ps@HP�s��?             9@�       �                   �`@�nkK�?             7@�       �                    �?�C��2(�?             &@�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?և���X�?             ,@�       �                   �_@�����H�?             "@�       �                   �r@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B0       �y@     �@     0t@     `o@     �H@     �j@      H@      c@      *@     �]@       @      ,@      �?              @      ,@      �?       @      �?      @      �?       @               @      �?                      @               @      @      @      @      @              @      @              @      @      �?      @      �?      �?              �?      �?                       @       @              @     @Z@       @     @Y@             �K@       @      G@       @      $@      �?              �?      $@      �?      @              @      �?                      @              B@      @      @               @      @       @               @      @             �A@     �@@      @      0@       @      @              @       @              �?      *@      �?                      *@      @@      1@      @@      *@      :@      @               @      :@       @      :@      �?      7@              @      �?      @                      �?              �?      @      "@      @      @      @              @      @      @                      @              @              @      �?     �O@      �?       @              @      �?      �?              �?      �?                     �K@      q@      B@      @      .@      @      @      @      �?              �?      @              �?      @      �?      �?              �?      �?                      @              $@     �p@      5@      D@      &@      D@      @      @      @      @              �?      @      �?       @               @      �?                      @     �@@      �?      .@      �?       @              @      �?      @      �?      @                      �?      @              2@                      @     �l@      $@      I@      @      F@      �?      =@              .@      �?              �?      .@              @      @      @      �?              �?      @                      @     �f@      @     �c@      �?     �E@             �\@      �?     �Q@      �?      Q@      �?      P@              @      �?      @                      �?       @              F@              7@       @      @       @               @      @              2@             �V@     �o@      ;@      @@      @      9@      @      "@               @      @      �?       @      �?       @                      �?      @                      0@      6@      @      �?      @      �?                      @      5@             �O@     �k@      :@     �f@      $@     @a@              B@      $@     �Y@      @      (@      @       @       @              @       @               @      @                      $@      @     �V@      @      B@      @      &@              "@      @       @       @              @       @              �?      @      �?       @              �?      �?      �?                      �?              9@              K@      0@      E@      @      @@      �?      5@      �?      @      �?                      @              .@      @      &@      @                      &@      &@      $@      "@      @              @      "@               @      @       @      �?       @                      �?              @     �B@      E@      �?      &@      �?       @      �?                       @              "@      B@      ?@      @      0@      @      @      @      @      @               @      @               @       @      �?      �?              �?      �?              �?      �?                       @              &@      ?@      .@      9@      @      7@       @      6@      �?      $@      �?      @      �?      @                      �?      @              (@              �?      �?      �?                      �?       @      @       @                      @      @       @      �?       @      �?       @      �?                       @              @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ\�0\hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK݅�h~�BX0         |       
             �?~jÚʞ�?Q           ��@       C                    �?<�A+K&�?O           ��@                           �?<�g���?�            �u@                          �a@�L"��?K            �Z@                          `_@z�G�z�?:            @U@       	                    �?ףp=
�?#             I@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?
                          Pr@=QcG��?             �G@������������������������       �                    �E@                          �\@      �?             @������������������������       �                     �?������������������������       �                     @                           �K@^������?            �A@                           �?��S�ۿ?	             .@������������������������       �                     �?������������������������       �                     ,@              	          ����?�G�z��?             4@������������������������       �                     @                           �?ҳ�wY;�?             1@                          �n@"pc�
�?             &@������������������������       �                     @                           �?      �?             @������������������������       �                      @������������������������       �                      @                          �w@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     6@       @                    �R@�U:�h�?�             n@        /                    j@P�H�}��?�            �m@!       .                    �L@���.�6�?@             W@"       #       	          033�?      �?"             H@������������������������       �                     8@$       '                    \@      �?             8@%       &                    g@      �?             @������������������������       �                     �?������������������������       �                     @(       -                    �?R���Q�?             4@)       ,       	          ����?d}h���?             ,@*       +                    �C@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     @������������������������       �                     F@0       ?       	          ��� @�-�|�?\            `b@1       >                   (q@����q�?E            @[@2       7                    �H@h㱪��?$            �K@3       6                    �?ףp=
�?             $@4       5                   �k@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @8       9                   �p@����?�?            �F@������������������������       �                     D@:       ;                   `a@z�G�z�?             @������������������������       �                     @<       =                   @^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        !             K@������������������������       �                     C@A       B                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?D       K                    �? �]^m>�?f             g@E       H                    �?ܷ��?��?             =@F       G                    @ �q�q�?             8@������������������������       �                     7@������������������������       �                     �?I       J                   �o@���Q��?             @������������������������       �                     @������������������������       �                      @L       m                   �b@��/W�?W            `c@M       N                   @Y@�S����?@            �\@������������������������       �                      @O       P                   �]@؇���X�??             \@������������������������       �                     :@Q       b                    �?&^�)b�?-            �U@R       S                   �\@�5��
J�?             G@������������������������       �                      @T       U       
             �?p9W��S�?             C@������������������������       �                     @V       Y                    �?H�V�e��?             A@W       X                   �c@�q�q�?             @������������������������       �                     @������������������������       �                      @Z       [                   0b@ �Cc}�?             <@������������������������       �                     2@\       _                    �?�z�G��?             $@]       ^                    @N@���Q��?             @������������������������       �                      @������������������������       �                     @`       a                   �`@z�G�z�?             @������������������������       �                     �?������������������������       �                     @c       d                    @M@      �?             D@������������������������       �                     8@e       f                    �?     ��?             0@������������������������       �                     @g       h                   @^@�q�q�?             (@������������������������       �                     @i       l                    `@      �?              @j       k                   �`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @n       o                   �c@�p ��?            �D@������������������������       �                     @p       {                    �?և���X�?            �A@q       x                   p@     ��?             @@r       u       	          ���@p�ݯ��?             3@s       t                   `e@r�q��?             (@������������������������       �                      @������������������������       �                     $@v       w                    �B@����X�?             @������������������������       �                      @������������������������       �                     @y       z                   f@�θ�?             *@������������������������       �                     $@������������������������       �                     @������������������������       �                     @}       �                    �?ʨ����?            x@~       �                    P@��+��?S            �[@       �                    �?��a�n`�?             ?@�       �                   �b@��s����?             5@�       �                     E@�8��8��?             (@�       �                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                   c@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �L@�z�G��?             $@������������������������       �                     @�       �                   @_@���Q��?             @�       �                    �?�q�q�?             @�       �                   �V@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    �?      �?>             T@�       �                    �D@�MWl��?+            �L@�       �                    @C@�eP*L��?             &@������������������������       �                     @�       �                   �b@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?�㙢�c�?$             G@�       �                    �?� ��1�?             �D@������������������������       �                     @�       �                   �a@4�2%ޑ�?            �A@�       �                   pa@�X�<ݺ?             2@������������������������       �        	             (@�       �                    �?r�q��?             @�       �                    `P@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �                    �?j���� �?             1@�       �                   pm@և���X�?             @������������������������       �                      @�       �       	          ����?z�G�z�?             @�       �                   p`@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   �_@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          ����?��+7��?             7@�       �                    b@X�<ݚ�?             "@������������������������       �                      @�       �                   (p@և���X�?             @�       �                    h@z�G�z�?             @������������������������       �                      @�       �                   �d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                   @_@@4և���?             ,@�       �                   �t@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �       	          ���@��Mj��?�            0q@�       �                    I@�ne�!2�?�            �p@�       �       	          ����?X�<ݚ�?             "@�       �                    `Q@r�q��?             @������������������������       �                     @�       �                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �L@�z�N��?�            `p@�       �                   �_@@p�<��?�             k@�       �                   @c@ �q�q�?             8@������������������������       �                     �?������������������������       �                     7@������������������������       �        t             h@�       �                     P@�q��/��?             G@�       �                    �?�חF�P�?             ?@�       �                    �O@�>4և��?             <@�       �                   `p@HP�s��?             9@������������������������       �                     2@�       �                   `c@����X�?             @�       �                    `@r�q��?             @������������������������       �                     @�       �                   �r@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        
             .@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       �y@     �@     �V@     �{@      :@      t@      1@     �V@      1@      Q@      @     �F@       @      �?       @                      �?      @      F@             �E@      @      �?              �?      @              (@      7@      �?      ,@      �?                      ,@      &@      "@              @      &@      @      "@       @      @               @       @       @                       @       @      @              @       @                      6@      "@      m@       @     �l@      @     �U@      @      E@              8@      @      2@      @      �?              �?      @              @      1@      @      &@      @      �?              �?      @                      $@              @              F@       @      b@       @     �Z@       @     �J@      �?      "@      �?      �?              �?      �?                       @      �?      F@              D@      �?      @              @      �?      �?              �?      �?                      K@              C@      �?      �?              �?      �?             @P@     �]@      :@      @      7@      �?      7@                      �?      @       @      @                       @     �C@      ]@      2@      X@       @              0@      X@              :@      0@     �Q@      &@     �A@               @      &@      ;@      @              @      ;@      @       @      @                       @      @      9@              2@      @      @       @      @       @                      @      �?      @      �?                      @      @     �A@              8@      @      &@              @      @      @      @              �?      @      �?       @               @      �?                      @      5@      4@      @              .@      4@      .@      1@      (@      @      $@       @               @      $@               @      @       @                      @      @      $@              $@      @                      @     �s@      Q@     �L@      K@      @      8@      @      1@      �?      &@      �?      �?              �?      �?                      $@      @      @              @      @              @      @              @      @       @      �?       @      �?      �?              �?      �?                      �?       @              I@      >@      F@      *@      @      @      @              �?      @      �?                      @      C@       @     �@@       @      @              ;@       @      1@      �?      (@              @      �?      @      �?      @                      �?       @              $@      @      @      @       @              �?      @      �?       @               @      �?                       @      @      @              @      @              @              @      1@      @      @       @              @      @      �?      @               @      �?       @               @      �?               @              �?      *@      �?      @              @      �?                       @     Pp@      ,@     Pp@      $@      @      @      @      �?      @              �?      �?      �?                      �?              @      p@      @     �j@      �?      7@      �?              �?      7@              h@             �D@      @      :@      @      7@      @      7@       @      2@              @       @      @      �?      @               @      �?       @                      �?              �?              @      @              .@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ+BhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B(5         �       
             �?z�ГPo�?1           ��@       +                    �?�:��a�??           ��@       *                    �?7�A�0�?4             V@       #                   �b@������?+            @Q@              	             �?�q�q�?              K@                          q@������?            �F@                           �?"pc�
�?            �@@       	                     L@ȵHPS!�?             :@������������������������       �        
             1@
                          k@�q�q�?             "@������������������������       �                     @                           �L@      �?             @������������������������       �                      @              	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?                          k@և���X�?             @������������������������       �                      @                          �]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                           �?      �?             (@������������������������       �                     @                           �?؇���X�?             @������������������������       �                     @                           �?      �?             @                          �r@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?                             K@�q�q�?             "@������������������������       �                      @!       "                    �O@؇���X�?             @������������������������       �                     @������������������������       �                     �?$       )       	             �?��S�ۿ?             .@%       (                   `c@�����H�?             "@&       '                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        	             3@,       �                   f@�wAf��?           �{@-       8       	          833�?8��8���?            {@.       /                    �K@�K}��?9            �Y@������������������������       �                    �I@0       7                    �?���J��?            �I@1       2                    �?��?^�k�?            �A@������������������������       �                     8@3       6                   @_@�C��2(�?             &@4       5                    @M@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �        
             0@9       v                    �?�r����?�            �t@:       M                    �?Hm_!'1�?�            �n@;       F                   pb@D>�Q�?             J@<       C                    `@������?            �D@=       >                   @^@���!pc�?             &@������������������������       �                      @?       @                   �]@�����H�?             "@������������������������       �                     @A       B                    �I@      �?              @������������������������       �                     �?������������������������       �                     �?D       E                   `x@(;L]n�?             >@������������������������       �                     =@������������������������       �                     �?G       L                    �?�eP*L��?             &@H       K                    �?����X�?             @I       J                   �r@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @N       O                   �U@�0p<���?z             h@������������������������       �                     �?P       U                    �?p�qG�?y             h@Q       T                   �Z@�Ń��̧?             E@R       S       	          033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     D@V       _                    \@ "��u�?a            �b@W       X                   ph@"pc�
�?             &@������������������������       �                     @Y       Z                   Pk@�q�q�?             @������������������������       �                     �?[       \                    �?z�G�z�?             @������������������������       �                     @]       ^       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?`       o                   �b@PX�V|�?Y            `a@a       f       	          033�?T��,��?A            @Y@b       e                    �?r�q��?             @c       d                    @J@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @g       j                   �X@ r���?>            �W@h       i                   �W@      �?             @������������������������       �                     @������������������������       �                     �?k       n                    _@@��,B�?:            �V@l       m                    \@$�q-�?
             *@������������������������       �                     �?������������������������       �        	             (@������������������������       �        0            �S@p       u                     R@�KM�]�?             C@q       t                   �f@�X�<ݺ?             B@r       s                   `U@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     ?@������������������������       �                      @w       �                   P`@Gq����?5            @U@x       �       	          033�?~�4_�g�?             F@y       z                   �Z@�ʻ����?             A@������������������������       �                     @{       |                   �k@l��
I��?             ;@������������������������       �                     ,@}       ~       
             �?�n_Y�K�?
             *@������������������������       �                      @       �                   �r@���!pc�?	             &@�       �                    �D@z�G�z�?             $@������������������������       �                     �?�       �                    �?�����H�?             "@������������������������       �                     @�       �                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                    �?,���i�?            �D@�       �                   �`@�z�G��?             $@������������������������       �                     @�       �       
             �?      �?             @������������������������       �                      @�       �                   c@      �?             @������������������������       �                     �?�       �                   `c@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   �T@`Jj��?             ?@�       �       	             �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     ;@�       �                   `e@������?             .@������������������������       �                     @�       �       	             @�8��8��?             (@������������������������       �                     &@������������������������       �                     �?�       �                    �?^��/O��?�            �w@�       �       	          ����?&ޑ���?Y            �a@�       �                    �?\`*�s�?5             U@�       �                    @F@�eP*L��?             6@������������������������       �                      @�       �                   �o@����X�?
             ,@������������������������       �                     @�       �                   �`@      �?              @�       �                    ^@�q�q�?             @������������������������       �                     �?�       �                   Pc@z�G�z�?             @������������������������       �                      @�       �                   �r@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �                    `@t�7��?)             O@�       �                   �[@R�}e�.�?             :@�       �                   @V@      �?              @������������������������       �                     �?�       �                   �Z@և���X�?             @�       �                    �J@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �_@r�q��?             2@�       �                   �Y@      �?             0@������������������������       �                     �?������������������������       �                     .@������������������������       �                      @�       �                   �c@�����H�?             B@������������������������       �                     8@�       �                    �?�q�q�?             (@�       �                   @d@z�G�z�?             $@������������������������       �                     �?�       �                    �?�����H�?             "@�       �                   @b@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   �u@d}h���?$             L@�       �                    X@�iʫ{�?"            �J@�       �                    _@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   0e@8��8���?              H@�       �                     P@��S�ۿ?            �F@�       �                    @K@������?             B@�       �                    �J@$�q-�?
             *@������������������������       �        	             (@������������������������       �                     �?������������������������       �                     7@�       �                    �?�<ݚ�?             "@�       �                   �m@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �V@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    I@ ��� �?�            `n@�       �                    �Q@���Q��?             @������������������������       �                     �?�       �                   �]@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �L@0x�!���?�            �m@�       �                   c@�K��h�?}            �h@�       �                   �b@�zvܰ?:             V@������������������������       �        9            @U@������������������������       �                     @������������������������       �        C            �[@�       �                   `b@�ݜ�?            �C@�       �                   �s@д>��C�?             =@�       �       	             �?$�q-�?             :@�       �                    d@`2U0*��?             9@������������������������       �                     2@�       �                    �?؇���X�?             @������������������������       �                     @�       �                     @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B0       �x@     @�@     @W@     �{@     �B@     �I@     �B@      @@      B@      2@     �@@      (@      ;@      @      7@      @      1@              @      @      @              �?      @               @      �?      �?      �?                      �?      @      @               @      @      �?              �?      @              @      @      @              �?      @              @      �?      @      �?       @               @      �?                      �?      @      @       @              �?      @              @      �?              �?      ,@      �?       @      �?      �?              �?      �?                      @              @              3@      L@     px@     �F@     0x@      �?     @Y@             �I@      �?      I@      �?      A@              8@      �?      $@      �?      @      �?                      @              @              0@      F@     �q@      4@      l@      "@     �E@      @     �B@      @       @       @              �?       @              @      �?      �?      �?                      �?      �?      =@              =@      �?              @      @      @       @      �?       @               @      �?              @                      @      &@     �f@      �?              $@     �f@      �?     �D@      �?      �?              �?      �?                      D@      "@     �a@       @      "@              @       @      @      �?              �?      @              @      �?      �?      �?                      �?      @     �`@      @     �X@      �?      @      �?       @               @      �?                      @       @     @W@      �?      @              @      �?              �?     �V@      �?      (@      �?                      (@             �S@      @      A@       @      A@       @      @              @       @                      ?@       @              8@     �N@      3@      9@      3@      .@              @      3@       @      ,@              @       @       @              @       @       @       @      �?              �?       @              @      �?       @               @      �?              �?                      $@      @      B@      @      @              @      @      @       @              �?      @              �?      �?       @               @      �?               @      =@       @       @       @                       @              ;@      &@      @              @      &@      �?      &@                      �?     s@     �S@     @R@     �P@     �N@      7@      $@      (@               @      $@      @      @              @      @       @      @      �?              �?      @               @      �?       @               @      �?               @             �I@      &@      3@      @      @      @      �?              @      @      �?      @      �?                      @       @              .@      @      .@      �?              �?      .@                       @      @@      @      8@               @      @       @       @              �?       @      �?      @      �?      @                      �?      @                       @      (@      F@      "@      F@      @      �?      @                      �?      @     �E@      @      E@      �?     �A@      �?      (@              (@      �?                      7@       @      @       @      @       @                      @              �?       @      �?              �?       @              @              m@      &@       @      @      �?              �?      @      �?                      @     �l@       @     �h@      @     @U@      @     @U@                      @     �[@              A@      @      8@      @      8@       @      8@      �?      2@              @      �?      @              @      �?      @                      �?              �?              @      $@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�vhkhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�<         �                    �?TU�`��?<           ��@       �                    �?t:ɨ2�?O           ��@       �       	          033�?�ͭ�1��?           py@       E                    �?��K��?�            �w@                          �_@���q��?R            �]@              
             �?��J�fj�?            �B@       
                    �?؇���X�?             5@       	                   �m@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     1@                           �J@     ��?             0@                          `]@�C��2(�?             &@������������������������       �                      @                          �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �M@���Q��?             @                          �X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @       D                   �{@�4F����?:            �T@       +       
             �?�J�j�?8            �S@       "                   �b@��
ц��?             :@                           X@�θ�?             *@������������������������       �                     �?              	          ����?r�q��?             (@������������������������       �                     �?                           b@�C��2(�?             &@������������������������       �                      @        !                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @#       *                   �e@�	j*D�?	             *@$       )                    �N@"pc�
�?             &@%       (                    o@ףp=
�?             $@&       '       	             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                      @,       -                    �? {��e�?'            �J@������������������������       �        	             ,@.       7                    ]@�(�Tw��?            �C@/       4                   �b@���Q��?             $@0       1                   �[@      �?             @������������������������       �                     �?2       3                   �a@�q�q�?             @������������������������       �                     �?������������������������       �                      @5       6                   �k@r�q��?             @������������������������       �                     �?������������������������       �                     @8       =                   d@д>��C�?             =@9       <                    �G@�}�+r��?             3@:       ;       	          ����?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             ,@>       C                   �b@���Q��?             $@?       @                   �^@      �?              @������������������������       �                     @A       B                   �l@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @F       S                    c@�s�,�?�            Pp@G       L                   �\@���Q��?             .@H       I                    @K@z�G�z�?             @������������������������       �                     @J       K                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?M       N                    �?z�G�z�?             $@������������������������       �                     �?O       R       	          ����?�����H�?             "@P       Q                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @T       w                    @L@���>�?�            �n@U       v                   �~@��'cy�?x            @i@V       c                    �?�/��5�?w             i@W       X                    �G@�h����?E             \@������������������������       �                     �L@Y       \                    @H@h㱪��?%            �K@Z       [                   �m@�q�q�?             @������������������������       �                     �?������������������������       �                      @]       ^                    �J@ pƵHP�?"             J@������������������������       �                     5@_       b                    �?�g�y��?             ?@`       a                   `f@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@d       q       	          ����?�ƫ�%�?2            @V@e       f                    @G@��pBI�?)            @R@������������������������       �                    �E@g       h                   �b@��S�ۿ?             >@������������������������       �        
             ,@i       j                    �?      �?             0@������������������������       �                     @k       p                    �?8�Z$���?             *@l       o                    o@z�G�z�?             $@m       n                   �^@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @r       u                    @     ��?	             0@s       t       	             �?�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     �?x       {                   �_@      �?             F@y       z                    �?      �?             @������������������������       �                     �?������������������������       �                     @|       �                   @t@z�G�z�?             D@}       �                    �?:�&���?            �C@~       �       
             �?���7�?             6@       �       	          pff�?�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     *@�       �       	          pff�?ҳ�wY;�?             1@�       �       	          @33�?r�q��?	             (@�       �                    @�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                     M@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �                    `P@X�<ݚ�?             ;@�       �                    �?����X�?             5@������������������������       �        	             *@�       �                   �a@      �?              @������������������������       �                     �?�       �                    �?؇���X�?             @�       �       	          `ff@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       
             �?*AA,�P�?L            @^@�       �                   �x@H%u��?/            �R@�       �                    �?�ӖF2��?.            �Q@�       �       
             �?      �?              @������������������������       �                      @������������������������       �                     @�       �                   �k@���N8�?*            �O@������������������������       �        !             G@�       �                   �n@@�0�!��?	             1@������������������������       �                     @������������������������       �                     ,@������������������������       �                     @�       �                    �?\X��t�?             G@�       �       	             �?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?�       �                    �?���@M^�?             ?@������������������������       �        	             ,@�       �                   ``@�t����?             1@������������������������       �                     @�       �                    �M@$�q-�?             *@������������������������       �        	             &@�       �                   `a@      �?              @������������������������       �                     �?������������������������       �                     �?�              
             �?L�B{�?�            `x@�       �                    �R@,��>��?�            �u@�       �                   pa@�{�{t��?�            Pu@�       �       	             �?xh�ڝ�?�            �p@������������������������       �        !            �J@�       �                    �?�V���?�            �j@�       �       	          ����?@�E�x�?W            `b@�       �                   �d@�nkK�?)            @Q@������������������������       �                     4@�       �                   �e@��<D�m�?            �H@������������������������       �                     �?�       �                    �? �q�q�?             H@�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?�       �                   @^@`���i��?             F@�       �                   �\@�C��2(�?             &@������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                    �@@������������������������       �        .            �S@�       �                   �`@l��\��?)             Q@�       �                    �?���B���?             :@�       �                    @J@�t����?	             1@������������������������       �                     @�       �                    r@�eP*L��?             &@�       �                    �?      �?              @������������������������       �                     �?�       �                    �J@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     "@�       �                   �u@�Ń��̧?             E@������������������������       �                     D@�       �                    @L@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�1��u�?,            @R@�       �                   �a@�X�C�?              L@�       �       	          hff�?���"͏�?            �B@�       �                    _@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �a@"pc�
�?            �@@�       �                    ^@      �?              @������������������������       �                     @�       �                   �f@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �Z@HP�s��?             9@������������������������       �                     �?�       �                    a@ �q�q�?             8@������������������������       �        	             3@�       �                   �n@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@�       �                   p@ҳ�wY;�?             1@�       �                    �?8�Z$���?             *@������������������������       �                     @�       �                    �E@z�G�z�?             $@������������������������       �                      @�       �                    �?      �?              @������������������������       �                      @�       �                    �?�q�q�?             @�       �                    �H@      �?             @������������������������       �                     �?�       �                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       	             @      �?             @������������������������       �                     @������������������������       �                     �?                         `@F�����?            �F@                        �W@      �?             0@������������������������       �                     �?                        �d@��S�ۿ?
             .@������������������������       �        	             ,@������������������������       �                     �?                        �j@l��[B��?             =@                         �?�t����?             1@	                         @N@�n_Y�K�?	             *@
                         �M@      �?              @                         a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @                         �?r�q��?             (@                        `@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�t�b�m7     h�h(h+K ��h-��R�(KMKK��h_�BP       @y@     �@     0v@     �e@      t@     �U@     @s@      R@      R@     �G@      0@      5@      @      2@      @      �?              �?      @                      1@      *@      @      $@      �?       @               @      �?              �?       @              @       @      �?       @               @      �?               @              L@      :@      L@      7@      ,@      (@      $@      @              �?      $@       @              �?      $@      �?       @               @      �?              �?       @              @      "@       @      "@      �?      "@      �?       @               @      �?                      @      �?               @              E@      &@      ,@              <@      &@      @      @      @      �?      �?               @      �?              �?       @              �?      @      �?                      @      8@      @      2@      �?      @      �?      @                      �?      ,@              @      @      @       @      @              @       @               @      @                       @              @     �m@      9@      "@      @      �?      @              @      �?      �?      �?                      �?       @       @              �?       @      �?       @      �?              �?       @              @             `l@      3@     @h@       @     @h@      @     �[@       @     �L@             �J@       @       @      �?              �?       @             �I@      �?      5@              >@      �?      @      �?      @                      �?      ;@              U@      @     �Q@       @     �E@              <@       @      ,@              ,@       @      @              &@       @       @       @      @       @               @      @              @              @              *@      @      @      @              @      @              @                      �?     �@@      &@      �?      @      �?                      @      @@       @      @@      @      5@      �?       @      �?       @                      �?      *@              &@      @      $@       @      @       @      @                       @      @              �?      @      �?                      @              �?      (@      .@      @      .@              *@      @       @              �?      @      �?      @      �?       @              �?      �?      �?                      �?      @              @             �A@     �U@      "@     �P@      @     �P@       @      @       @                      @      @      N@              G@      @      ,@      @                      ,@      @              :@      4@      ,@      �?      ,@                      �?      (@      3@              ,@      (@      @              @      (@      �?      &@              �?      �?      �?                      �?     �H@     Pu@      @@     �s@      =@     �s@      "@     0p@             �J@      "@     �i@      @      b@      @     �P@              4@      @      G@      �?               @      G@      �?      @              @      �?              �?     �E@      �?      $@               @      �?       @      �?                       @             �@@             �S@      @      O@      @      5@      @      (@              @      @      @       @      @              �?       @      @       @                      @      @                      "@      �?     �D@              D@      �?      �?              �?      �?              4@     �J@      "@     �G@      "@      <@      @      �?              �?      @              @      ;@      @      @      @              �?      @      �?                      @       @      7@      �?              �?      7@              3@      �?      @              @      �?                      3@      &@      @      &@       @      @               @       @       @              @       @       @              @       @       @       @              �?       @      �?       @                      �?       @                      @      @      �?      @                      �?      1@      <@       @      ,@      �?              �?      ,@              ,@      �?              .@      ,@      @      (@      @       @      @      @      �?      @      �?                      @      @                      @              @      $@       @       @       @       @                       @       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJF�3hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM1hwh(h+K ��h-��R�(KM1��h~�B�B         �       
             �?�$�����?P           ��@       M                   P`@ %团��?T           �@       F                    �?(�7T�<�?�            �r@       1                   P`@8Fb����?�            @i@                           `@6�����?H            @[@                           �?�F��O�?3            @R@                           ]@���Q��?             @������������������������       �                      @	       
                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @                           �? =[y��?.             Q@                           �?�KM�]�?             3@                          �]@�X�<ݺ?             2@������������������������       �                     @                          �W@$�q-�?             *@                           �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?              	          033@@�E�x�?"            �H@������������������������       �                     E@                          �^@؇���X�?             @������������������������       �                     @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?       $                    @L@�q�q�?             B@       #                    ^@      �?             0@                            �?      �?              @������������������������       �                     �?!       "       	          033�?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @%       &                    �?�G�z��?
             4@������������������������       �                      @'       ,                    �?b�2�tk�?	             2@(       )                    [@����X�?             @������������������������       �                     �?*       +                   �^@r�q��?             @������������������������       �                     @������������������������       �                     �?-       0                   `]@�eP*L��?             &@.       /                    �L@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @2       E                   �b@�g�y��?A            @W@3       8                    �D@���N8�?.            �O@4       7       	             �?�q�q�?             @5       6                    �C@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?9       >                    �?(;L]n�?+             N@:       ;                    �?      �?             @������������������������       �                     �?<       =                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �??       D                   �a@�h����?(             L@@       C                    @L@Pa�	�?            �@@A       B       	          ����?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     5@������������������������       �                     7@������������������������       �                     >@G       L       	          ����?�����?@            @Y@H       K       
             �? �Jj�G�?#            �K@I       J                   �l@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        !            �J@������������������������       �                     G@N       �                    �?#z�i��?�            �i@O       ~                   �b@���hg��?c            �b@P       {       	          `ff@DrfuN�?>            �W@Q       j                    �?���!pc�?<             V@R       U       
             �?r�q��?(             N@S       T       	             @z�G�z�?             $@������������������������       �                      @������������������������       �                      @V       a                    �?�J�4�?"             I@W       `                   �p@���|���?	             &@X       Y                   �`@և���X�?             @������������������������       �                      @Z       _                   �o@���Q��?             @[       ^                   �g@      �?             @\       ]                     M@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @b       e                    @I@��-�=��?            �C@c       d                    �F@�z�G��?             $@������������������������       �                     @������������������������       �                     @f       i                   h@XB���?             =@g       h       	          ����?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     7@k       r                   0l@      �?             <@l       q                    �?r�q��?	             (@m       n       	          833�?����X�?             @������������������������       �                     @o       p                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @s       x                    �M@      �?             0@t       u       	          @33�?8�Z$���?	             *@������������������������       �                     @v       w                    �?      �?              @������������������������       �                      @������������������������       �                     @y       z                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?|       }                    e@r�q��?             @������������������������       �                     �?������������������������       �                     @       �                   c@X�<ݚ�?%             K@������������������������       �                     $@�       �                   �f@�eP*L��?             F@�       �                   p@���Q��?             D@�       �                    �?|��?���?             ;@�       �                    �?      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?�       �       	          `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �K@p�ݯ��?             3@�       �       	          ����?r�q��?	             (@������������������������       �                     @�       �                   �d@���Q��?             @������������������������       �                      @������������������������       �                     @�       �                   �c@����X�?             @�       �                     O@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?�θ�?
             *@�       �       	          ���@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?�����H�?             "@������������������������       �                     @�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     Q@F�t�K��?(            �L@�       �                    �?�2����?'            �K@�       �                    �K@��?^�k�?            �A@������������������������       �                     1@�       �                    �?�X�<ݺ?             2@������������������������       �                     ,@�       �                     M@      �?             @������������������������       �                     �?������������������������       �                     @�       �                   �a@���Q��?             4@�       �                   `_@������?             .@�       �       
             �?      �?             @������������������������       �                     �?�       �       	          ����?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �c@�����H�?             "@�       �                    �?      �?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �d@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�                          �?� ��1�?�            �y@�       �                    @K@�ʻ����?Q             a@�       �                    f@�	j*D�?-            �S@�       �                   �_@����X�?	             ,@�       �                   @[@r�q��?             (@�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       �                   �b@     ��?$             P@�       �                   �a@��S�ۿ?             >@�       �                    @G@ 7���B�?             ;@�       �       	          ����?�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     2@�       �                    �?�q�q�?             @������������������������       �                     �?�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �f@ҳ�wY;�?             A@�       �                    �?�q�����?             9@������������������������       �                     @�       �                    �?�eP*L��?             6@�       �                    �?      �?             4@������������������������       �                     @�       �                   �[@j���� �?             1@������������������������       �                     @�       �                   Pm@��
ц��?
             *@������������������������       �                     @�       �                   d@�q�q�?             "@������������������������       �                     @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     "@�                          �?����"�?$             M@�       �                   `a@
;&����?             G@�       �                   @E@$��m��?             :@�       �                    �?r�q��?             @�       �                    �?      �?             @������������������������       �                     �?�       �                   �X@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�       �       	          ����?z�G�z�?             4@�       �       	          ����?����X�?
             ,@�       �                    �?�C��2(�?             &@������������������������       �                     @�       �                    �L@      �?              @������������������������       �                     @�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �M@      �?             4@�       �                    �?և���X�?             @������������������������       �                     @�       �                    @M@      �?             @������������������������       �                     @������������������������       �                     �?�                           S@$�q-�?             *@�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@������������������������       �                     (@      .                  0h@ȥ�fzR�?�             q@                         �?��j���?�            �p@            	          833@�q��/��?            �H@                        �`@8��8���?             H@������������������������       �                    �@@      	                   �?�q�q�?             .@������������������������       �                     @
                         @M@r�q��?             (@������������������������       �                     @                          O@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?      '                   �?@-�_ .�?�            �k@      &                  Pd@��ɉ�?            `h@            	            �?���7�?T            �`@                         I@PԱ�l�?D            �Z@                        �b@z�G�z�?             $@������������������������       �                      @������������������������       �                      @                        �b@`�E���?>            @X@������������������������       �        .            @Q@                        @[@@4և���?             <@                         �H@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     8@                         �?HP�s��?             9@������������������������       �                     "@       !                  `a@      �?	             0@������������������������       �                     "@"      %                  �p@����X�?             @#      $                  �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �        +            �O@(      +                   �?�<ݚ�?             ;@)      *                  �O@�㙢�c�?             7@������������������������       �                     @������������������������       �                     3@,      -                  P`@      �?             @������������������������       �                      @������������������������       �                      @/      0                   d@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KM1KK��h_�B       `z@      @      W@      z@      6@     �q@      5@     �f@      2@     �V@      @     �P@      @       @       @              �?       @      �?                       @      @     @P@       @      1@      �?      1@              @      �?      (@      �?      @              @      �?                       @      �?              �?      H@              E@      �?      @              @      �?       @               @      �?              (@      8@      �?      .@      �?      @              �?      �?      @      �?                      @               @      &@      "@               @      &@      @      @       @              �?      @      �?      @                      �?      @      @       @      @       @                      @      @              @     �V@      @      N@      �?       @      �?      �?              �?      �?                      �?       @      M@      �?      @              �?      �?       @               @      �?              �?     �K@      �?      @@      �?      &@      �?                      &@              5@              7@              >@      �?      Y@      �?      K@      �?      �?              �?      �?                     �J@              G@     �Q@     �`@     �M@     @V@      =@     @P@      8@      P@      $@      I@       @       @       @                       @       @      E@      @      @      @      @       @               @      @      �?      @      �?      �?      �?                      �?               @      �?                      @      @     �A@      @      @              @      @              �?      <@      �?      @              @      �?                      7@      ,@      ,@      $@       @      @       @      @              �?       @      �?                       @      @              @      (@       @      &@              @       @      @       @                      @       @      �?       @                      �?      @      �?              �?      @              >@      8@      $@              4@      8@      0@      8@      *@      ,@      @       @      �?       @              �?      �?      �?              �?      �?              @              @      (@       @      $@              @       @      @       @                      @      @       @      �?       @               @      �?              @              @      $@       @       @       @                       @      �?       @              @      �?      �?              �?      �?              @              &@      G@      "@      G@      �?      A@              1@      �?      1@              ,@      �?      @      �?                      @       @      (@      @      &@      @      @      �?               @      @              @       @              �?       @      �?      @      �?      �?      �?                      �?               @              @      @      �?      @                      �?       @             �t@      T@      S@      N@      K@      8@      @      $@       @      $@       @       @       @                       @               @       @              I@      ,@      <@       @      :@      �?       @      �?       @                      �?      2@               @      �?      �?              �?      �?      �?                      �?      6@      (@      *@      (@      @              $@      (@      $@      $@              @      $@      @      @              @      @              @      @      @      @              @      @      @                      @               @      "@              6@      B@      6@      8@      1@      "@      �?      @      �?      @              �?      �?       @               @      �?                       @      0@      @      $@      @      $@      �?      @              @      �?      @               @      �?       @                      �?              @      @              @      .@      @      @      @              �?      @              @      �?              �?      (@      �?      �?      �?                      �?              &@              (@     �o@      4@     �o@      2@     �E@      @     �E@      @     �@@              $@      @              @      $@       @      @              @       @               @      @                      �?     @j@      (@     �g@      @     �_@      @     �Y@      @       @       @       @                       @     �W@       @     @Q@              :@       @       @       @               @       @              8@              7@       @      "@              ,@       @      "@              @       @      �?       @      �?                       @      @             �O@              5@      @      3@      @              @      3@               @       @       @                       @      �?       @      �?                       @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ:%hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�9         �       
             �?������?1           ��@       i                   �b@@y��K��?G           ��@              	          ����?0=Aw�?           p{@                           �?@uvI��?<            �X@������������������������       �        )            �Q@                           �?h�����?             <@       
                    �H@؇���X�?             @       	                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     5@       F                   P`@"pc�
�?�            Pu@              	          ����?�Y��$�?�            �l@                          �[@�q�q�?             .@������������������������       �                      @                          �p@�θ�?             *@                           �?�C��2(�?             &@������������������������       �                     @              	          hff�?z�G�z�?             @                           @N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @       C                    �R@��hq��?�            �j@       B       	          pff�?|)���?�            @j@       ?                    �?x���� �?N             ^@              	          ����?z�G�z�?7             T@������������������������       �                      @       0                   �j@:�&���?5            �S@        !                    �?<ݚ)�?             B@������������������������       �                     @"       '       	          033�?r�q��?             >@#       &                   p`@�X�<ݺ?             2@$       %                   �X@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@(       -                    @L@�q�q�?             (@)       *                   �c@      �?              @������������������������       �                     @+       ,                    �C@�q�q�?             @������������������������       �                      @������������������������       �                     �?.       /                    �?      �?             @������������������������       �                     �?������������������������       �                     @1       >                    �?@4և���?             E@2       9                   @^@�#-���?            �A@3       8       	          ����? ��WV�?             :@4       7                    \@ףp=
�?	             $@5       6                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     0@:       ;                   �^@�<ݚ�?             "@������������������������       �                     �?<       =                    b@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @@       A                   �x@�(\����?             D@������������������������       �                    �C@������������������������       �                     �?������������������������       �        8            �V@D       E                   `c@      �?             @������������������������       �                     �?������������������������       �                     @G       \                    �?����X�?C             \@H       [                   ``@:�&���?+            �S@I       N                    �?p�ݯ��?             C@J       K                    @E@      �?              @������������������������       �                     �?L       M                    b@؇���X�?             @������������������������       �                     @������������������������       �                     �?O       R                   �j@������?             >@P       Q                   `[@�q�q�?             (@������������������������       �                     @������������������������       �                     @S       T                    �?r�q��?             2@������������������������       �                     @U       V                   �`@      �?             (@������������������������       �                      @W       Z                    \@ףp=
�?             $@X       Y                   �n@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     D@]       ^                    �?��.k���?             A@������������������������       �                     @_       `       
             �?և���X�?             <@������������������������       �                     @a       f                   b@��H�}�?             9@b       e                   �n@�n_Y�K�?
             *@c       d                     I@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                     @g       h                    _@�8��8��?	             (@������������������������       �                     �?������������������������       �                     &@j       �                    �? ��*��?7            �W@k       ~                   `a@���Q��?(            @P@l       u                   p@�	j*D�?             J@m       p                    @C@@�0�!��?             A@n       o                   pm@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @q       r                    @K@HP�s��?             9@������������������������       �                     2@s       t                    X@����X�?             @������������������������       �                      @������������������������       �                     @v       }                   �r@X�<ݚ�?             2@w       x                     G@�C��2(�?             &@������������������������       �                     @y       |                    �J@      �?             @z       {                   �p@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @       �                    �O@�θ�?	             *@�       �                    @G@�C��2(�?             &@�       �                   �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                      @�       �       	          ����?V�a�� �?             =@������������������������       �                     1@�       �                    �?      �?             (@������������������������       �                     @�       �                   �`@�q�q�?             "@�       �                   �X@؇���X�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �L@��K�R��?�            x@�       �                    �? U��?�            �q@�       �                   ``@�	j*D�?2            �S@�       �                   @E@�E��
��?             J@�       �                   `\@8�Z$���?             *@�       �       	             ��q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@�       �                   0o@��Sݭg�?            �C@�       �                   �a@�q�q�?             ;@������������������������       �                     &@�       �                   Pl@     ��?
             0@�       �       	             �?�q�q�?             "@�       �                    �C@և���X�?             @������������������������       �                      @�       �                    f@���Q��?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     �?�       �                    �G@�q�q�?             @������������������������       �                     �?�       �                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �l@؇���X�?             @������������������������       �                     @�       �       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �B@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�       �                   �c@ȵHPS!�?             :@�       �                    a@HP�s��?             9@������������������������       �                     $@�       �                    �K@�r����?             .@�       �                    @I@@4և���?             ,@������������������������       �                     @�       �                   �a@؇���X�?             @�       �       	          pff�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   �P@�g�A�E�?w            �i@�       �       	          ����?      �?              @������������������������       �                     @������������������������       �                     @�       �                    �?��:x�ٳ?t            �h@�       �                    c@r�q��?             8@�       �       	          pff�?���N8�?             5@������������������������       �                     1@�       �                   f@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    _@�d���?a            �e@�       �                   Hp@�kb97�?+            @S@������������������������       �        "             M@�       �                    �?���y4F�?	             3@������������������������       �                     &@�       �                    @K@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �        6            @X@�       �                    �?��H���?A            @Y@�       �                   @a@      �?             8@�       �                    �?      �?	             (@�       �                    �?      �?              @�       �                   a@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �        	             (@�       �       	          ����?��j��?/            @S@�       �                   hp@�4F����?            �D@�       �                    �?     ��?             @@�       �       	            �?�z�G��?             $@�       �                    �?�<ݚ�?             "@�       �                   �b@      �?              @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@�       �       	          @33�?�q�q�?             "@�       �                   �b@      �?              @�       �                   @c@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    `@r�q��?             B@������������������������       �        	             4@�                          �?      �?             0@�                          �?�eP*L��?             &@�              	          033	@X�<ݚ�?             "@�       �                    �?����X�?             @������������������������       �                      @�       �                    �?���Q��?             @�       �                    �M@      �?             @������������������������       �                     �?�       �       	          033�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                         @M@z�G�z�?             @������������������������       �                      @                         j@�q�q�?             @������������������������       �                      @������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KMKK��h_�Bp       �y@     �@      [@     �z@     �O@     �w@      �?     @X@             �Q@      �?      ;@      �?      @      �?      �?      �?                      �?              @              5@      O@     pq@      >@     �h@      $@      @               @      $@      @      $@      �?      @              @      �?      �?      �?              �?      �?              @                       @      4@     @h@      1@      h@      1@     �Y@      0@      P@       @              ,@      P@      &@      9@      @              @      9@      �?      1@      �?      @      �?                      @              $@      @       @      �?      @              @      �?       @               @      �?              @      �?              �?      @              @     �C@      @      @@      �?      9@      �?      "@      �?      @      �?                      @              @              0@       @      @      �?              �?      @              @      �?                      @      �?     �C@             �C@      �?                     �V@      @      �?              �?      @              @@      T@      ,@      P@      ,@      8@      @       @              �?      @      �?      @                      �?       @      6@      @      @      @                      @      @      .@              @      @      "@       @              �?      "@      �?      @      �?                      @              @              D@      2@      0@      @              (@      0@      @              "@      0@       @      @       @      �?              �?       @                      @      �?      &@      �?                      &@     �F@     �H@     �C@      :@      B@      0@      <@      @      @      @              @      @              7@       @      2@              @       @               @      @               @      $@      �?      $@              @      �?      @      �?      �?              �?      �?                       @      @              @      $@      �?      $@      �?      �?              �?      �?                      "@       @              @      7@              1@      @      @              @      @      @      @      �?      �?      �?              �?      �?              @                       @     �r@     �T@     �n@     �B@      K@      8@      ?@      5@       @      &@       @      �?              �?       @                      $@      =@      $@      2@      "@      &@              @      "@      @      @      @      @       @               @      @              �?       @       @              �?       @      �?      �?              �?      �?              �?      �?               @              �?      @              @      �?       @      �?                       @      &@      �?              �?      &@              7@      @      7@       @      $@              *@       @      *@      �?      @              @      �?       @      �?       @                      �?      @                      �?              �?      h@      *@      @      @      @                      @     �g@       @      4@      @      4@      �?      1@              @      �?              �?      @                      @     @e@      @     @R@      @      M@              .@      @      &@              @      @      @                      @     @X@             �K@      G@      5@      @      "@      @      @      @       @      @       @                      @      @              @              (@              A@     �E@      <@      *@      9@      @      @      @       @      @      �?      @      �?      �?      �?                      �?              @      �?              �?              6@              @      @       @      @       @       @       @                       @              @      �?              @      >@              4@      @      $@      @      @      @      @      @       @       @              @       @       @       @      �?              �?       @               @      �?              �?                       @               @      �?      @               @      �?       @               @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJr��hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B6         (                   �a@�&���?H           ��@              
             �?�[a���?z            �g@              	          033�? ��ʻ��?V             a@������������������������       �        :            �V@                          �c@`Ӹ����?            �F@������������������������       �                    �C@                           �?�q�q�?             @������������������������       �                     @	       
                   �d@�q�q�?             @������������������������       �                     �?                            M@      �?              @������������������������       �                     �?������������������������       �                     �?                          `@�1�`jg�?$            �K@              	          ����?�>����?             ;@                           �?����X�?             @������������������������       �                     @                          `[@      �?             @������������������������       �                     �?                          �`@�q�q�?             @������������������������       �                     �?                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     4@                          `a@      �?             <@                          �\@�8��8��?             (@                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@        '                   @E@     ��?             0@!       "                   �Y@�r����?
             .@������������������������       �                     �?#       $                   �b@@4և���?	             ,@������������������������       �                      @%       &                    �L@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?)       �                    �?��U����?�           ��@*       �                    �?��t�?�            �@+       d       
             �?��a^���?            `y@,       U                   `a@�w%�ob�?U             a@-       <                    �?�eP*L��?;             V@.       /       	          ����?�G�z�?             D@������������������������       �                     0@0       1                   �]@r�q��?             8@������������������������       �                     @2       3                    �?��Q��?             4@������������������������       �                     @4       7                   �]@��S���?
             .@5       6                   d@r�q��?             @������������������������       �                     @������������������������       �                     �?8       9                   �^@�<ݚ�?             "@������������������������       �                     @:       ;       	             �?���Q��?             @������������������������       �                     @������������������������       �                      @=       T                   d@r�qG�?              H@>       S                    �?�P�*�?             ?@?       D                    �?X�Cc�?             <@@       C                    �?ףp=
�?             $@A       B                    @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @E       F                   �e@      �?             2@������������������������       �                     @G       H                   l@���Q��?
             .@������������������������       �                     @I       R                   Pp@�q�q�?             "@J       K       	          ����?      �?             @������������������������       �                     �?L       Q                   �n@���Q��?             @M       N                    �?�q�q�?             @������������������������       �                     �?O       P                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     1@V       _                    @���c�H�?            �H@W       X                   �b@ףp=
�?             D@������������������������       �                     9@Y       Z                   0c@������?	             .@������������������������       �                     @[       \                   xu@�8��8��?             (@������������������������       �                     "@]       ^                   pc@�q�q�?             @������������������������       �                      @������������������������       �                     �?`       a                    �?�<ݚ�?             "@������������������������       �                     @b       c       
             �?      �?             @������������������������       �                      @������������������������       �                      @e       f                    �?����J��?�            �p@������������������������       �        :            �U@g       �                   �g@���'\�?q            �f@h       s                   �\@�����D�?p            �f@i       r                   m@��s����?             5@j       k                   @Z@���Q��?             $@������������������������       �                     @l       q                    �?և���X�?             @m       n                    �?z�G�z�?             @������������������������       �                     @o       p                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@t       �                   �t@      �?b             d@u       �                    �?=0�_�?_             c@v       }                    �?�S����?             3@w       |                   �q@����X�?             @x       {                   @p@r�q��?             @y       z                   �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?~                          @c@�8��8��?
             (@������������������������       �        	             &@������������������������       �                     �?�       �                    @5�wAd�?Q            �`@�       �                    @L@0�ޤ��?O            @`@�       �       	          ����? �O�H�?D            �[@������������������������       �        ?             Y@�       �                   �d@�C��2(�?             &@������������������������       �                     "@�       �       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �L@�KM�]�?             3@������������������������       �                      @������������������������       �        
             1@�       �                   �b@      �?             @������������������������       �                      @������������������������       �                      @�       �       	             �?����X�?             @�       �                    �J@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                   �c@Hя8X8�?�            �i@�       �                    �?�S1�<�?u            �g@�       �                    @G@�F���H�?g             e@�       �                   @n@�q�q�?             8@�       �                   �i@և���X�?	             ,@�       �                   �f@r�q��?             @�       �                   @e@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �`@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@�       �                   `\@      �?V             b@�       �                   `[@��0{9�?            �G@�       �                   �`@�g�y��?             ?@�       �                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �                     1@�       �       	          ����?      �?             0@������������������������       �                     @�       �                    �?r�q��?	             (@������������������������       �                     �?�       �                   Pn@�C��2(�?             &@������������������������       �                     @�       �                   �`@      �?             @������������������������       �                     �?������������������������       �                     @�       �       	          ����?`�E���?8            @X@�       �                    �?@9G��?            �H@�       �                    `@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   �i@�(\����?             D@�       �                   i@��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?������������������������       �                     9@������������������������       �                     H@�       �                   �[@���!pc�?             6@������������������������       �                     @�       �                   �b@�S����?             3@�       �       	          ����?�����H�?             2@�       �                    �K@      �?              @������������������������       �                     @�       �                   @_@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@������������������������       �                     �?�       �                   @l@      �?             0@�       �       	             �?ףp=
�?             $@�       �                     M@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    ]@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �       	          ����?�ʹ��Q�?M            �\@�       �                   �f@(옄��?!             G@������������������������       �                     @�       �       
             �?��
ц��?            �C@������������������������       �                     3@�       �                   �b@ףp=
�?             4@������������������������       �                     $@�       �                     I@z�G�z�?	             $@�       �                   �_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �J@��X���?,            @Q@�       �                    @H@��
ц��?
             *@������������������������       �                      @�       �                    d@���|���?             &@�       �                   P`@և���X�?             @�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       
             �? �Cc}�?"             L@�       �                    �L@�NW���?            �J@������������������������       �                     7@�       �                   �`@�r����?             >@������������������������       �                     �?�       �                   �l@ܷ��?��?             =@������������������������       �                     .@�       �                   pn@d}h���?             ,@������������������������       �                     @������������������������       �        	             &@�       �                   �`@�q�q�?             @������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�Bp        y@      �@      2@     �e@       @     �`@             �V@       @     �E@             �C@       @      @              @       @      �?      �?              �?      �?              �?      �?              0@     �C@       @      9@       @      @              @       @       @      �?              �?       @              �?      �?      �?              �?      �?                      4@      ,@      ,@      &@      �?      �?      �?      �?                      �?      $@              @      *@       @      *@      �?              �?      *@               @      �?      @              @      �?              �?              x@     pu@     �u@     �p@     �s@     @W@     �M@     �S@      H@      D@      *@      ;@              0@      *@      &@              @      *@      @      @               @      @      �?      @              @      �?              @       @      @              @       @      @                       @     �A@      *@      2@      *@      2@      $@      "@      �?      �?      �?      �?                      �?       @              "@      "@              @      "@      @      @              @      @      @      @              �?      @       @      �?       @              �?      �?      �?              �?      �?               @                      @              @      1@              &@      C@      @      B@              9@      @      &@      @              �?      &@              "@      �?       @               @      �?              @       @      @               @       @       @                       @     �o@      .@     �U@             �d@      .@     �d@      ,@      1@      @      @      @      @              @      @      �?      @              @      �?      �?      �?                      �?       @              &@             �b@      $@      b@       @      0@      @      @       @      @      �?       @      �?       @                      �?      @                      �?      &@      �?      &@                      �?      `@      @     �_@      @     �[@      �?      Y@              $@      �?      "@              �?      �?              �?      �?              1@       @               @      1@               @       @       @                       @      @       @       @       @       @                       @      @                      �?     �@@     �e@      7@     �d@      1@     �b@       @      0@       @      @      �?      @      �?      �?              �?      �?                      @      @      �?              �?      @                      $@      "@     �`@      @      D@      �?      >@      �?      *@              *@      �?                      1@      @      $@      @               @      $@      �?              �?      $@              @      �?      @      �?                      @       @     �W@       @     �G@      �?       @      �?                       @      �?     �C@      �?      ,@              ,@      �?                      9@              H@      @      0@      @              @      0@       @      0@       @      @              @       @      @              @       @                      $@      �?              $@      @      "@      �?      @      �?       @              �?      �?              �?      �?              @              �?      @      �?                      @      C@     @S@      9@      5@      @              2@      5@              3@      2@       @      $@               @       @       @       @       @                       @      @              *@      L@      @      @               @      @      @      @      @      @      �?      @                      �?              @      @              @      I@      @     �H@              7@      @      :@      �?              @      :@              .@      @      &@      @                      &@       @      �?              �?       @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJϩ�@hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B(<         <                    �?�O(�.��?V           ��@       -                    �?.��<�?x             i@                           @L@��}���?]            @c@                           �?����??            @Z@       
       	          ����?��8�$>�?;            @X@                          `c@�E�����?7            �V@������������������������       �        2            �T@       	                   �c@      �?              @������������������������       �                     �?������������������������       �                     @                           �?և���X�?             @                          Xq@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           @I@      �?              @                          �_@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @       "                   0c@ \� ���?            �H@                          �s@�ݜ�?            �C@                           �?�FVQ&�?            �@@              	          `ff @z�G�z�?             $@                          �e@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@       !                     P@      �?             @                           pc@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @#       ,                   0d@�z�G��?             $@$       %       
             �?�<ݚ�?             "@������������������������       �                     @&       '                   �c@�q�q�?             @������������������������       �                     �?(       +                    o@z�G�z�?             @)       *                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?.       7                   pn@"Ae���?            �G@/       0                    `@�q�q�?             2@������������������������       �                     @1       2                   �_@z�G�z�?	             .@������������������������       �                     �?3       6                    �?؇���X�?             ,@4       5                    V@$�q-�?             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?8       ;       	          ����?\-��p�?             =@9       :                   �[@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     8@=       �       
             �?��ė�X�?�           h�@>       a                   �g@4���t��?            �z@?       T                   Pe@����Q8�?g            �a@@       C                   �U@������?X            �^@A       B                    D@      �?              @������������������������       �                     �?������������������������       �                     �?D       Q                    �Q@���tcH�?V            @^@E       F                    �?���<_�?T            �]@������������������������       �        <            �U@G       N                    �?     ��?             @@H       M                   �`@8�Z$���?             *@I       J                   �Z@���Q��?             @������������������������       �                     �?K       L       	          `ff@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @O       P                   �e@�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?R       S                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?U       `                    c@�KM�]�?             3@V       _       	             �?؇���X�?             ,@W       ^                    �F@�<ݚ�?             "@X       Y                    �C@      �?             @������������������������       �                     �?Z       [                   �e@�q�q�?             @������������������������       �                     �?\       ]                   pf@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @b       �                    �?�HX���?�            �q@c       h       	          ����?f���M�?<            @W@d       g                   �i@�t����?             1@e       f                   �^@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@i       z                    �?��=A��?/             S@j       y                   �a@���?            �D@k       v                   (r@J�8���?             =@l       u                    �?��<b���?             7@m       t                   0a@"pc�
�?             6@n       o                    _@ףp=
�?             4@������������������������       �                      @p       s       	          ����?r�q��?             (@q       r                   0o@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     �?w       x       	          pff@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     (@{       �                   pf@���Q��?            �A@|       }       
             �?`՟�G��?             ?@������������������������       �                     @~                           �E@|��?���?             ;@������������������������       �                     @�       �                   Pp@�q�q�?             8@�       �       	            �?j���� �?	             1@������������������������       �                     @�       �                    �?�q�q�?             (@�       �                    �?      �?              @������������������������       �                     @�       �                    m@      �?             @������������������������       �                      @������������������������       �                      @�       �       	          pff@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                   �Z@X��R9�?}             h@�       �                   a@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?xrg��?z            �g@������������������������       �                     >@�       �                   0i@D���D|�?f            �c@�       �                   @`@�q�q�?             "@������������������������       �                     @������������������������       �                     @�       �                    �?Х-��ٹ?_            �b@�       �       
             �?�-�[�?Q            ``@�       �                   �\@�C��2(�?             6@�       �       	             �?�q�q�?             @������������������������       �                      @�       �                   �[@      �?             @������������������������       �                     �?�       �                   �c@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        	             0@�       �                    �M@��Ujѡ�?C            @[@�       �                   8q@@4և���?3             U@�       �                    c@lGts��?            �K@�       �                   �_@HP�s��?             I@�       �                   �^@z�G�z�?             .@�       �                   `a@�C��2(�?             &@������������������������       �                     @�       �                   �k@      �?             @������������������������       �                     @������������������������       �                     �?�       �       	             @      �?             @������������������������       �                      @������������������������       �                      @�       �                    @K@��?^�k�?            �A@������������������������       �                     7@�       �                   �a@�8��8��?             (@�       �       	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@�       �                   `c@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     =@������������������������       �                     9@������������������������       �                     3@�       �                   @E@�}*����?�            r@�       �       	          hff�?���Q��?             D@�       �                    �?�û��|�?             7@�       �                    �?"pc�
�?	             &@�       �                   �Y@      �?             @������������������������       �                     �?�       �                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       �                   c@�t����?             1@�       �       	          ����?      �?
             0@������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�                          �?�P{6�I�?�             o@�       �                    @L@�Z��L��?�            �j@�       �                    �?�y��`�?m            �e@�       �                    @J@��k=.��?            �G@�       �                    �I@��R[s�?            �A@�       �                    �?     ��?             @@�       �                   @^@      �?              @�       �       	          ����?z�G�z�?             @�       �                   `\@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �D@�8��8��?             8@�       �                    �C@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �                     0@������������������������       �                     @������������������������       �                     (@�       �                   @c@H�Swe�?O            @_@�       �                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                   �g@(;L]n�?L             ^@�       �                    �?@��,*�?K            �]@������������������������       �        ,            @Q@�       �                   @c@ "��u�?             I@�       �                    �G@؇���X�?             5@�       �                    @G@���!pc�?             &@������������������������       �                     @�       �                   �b@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     $@������������������������       �                     =@������������������������       �                     �?�                          �?��P���?            �D@�                         p@     ��?             @@�       �                    b@�LQ�1	�?             7@�       �       	          ����?@4և���?             ,@������������������������       �        
             *@������������������������       �                     �?�                          �?�<ݚ�?             "@�              	          `ff�?      �?             @�       �                    �?�q�q�?             @�       �                    �O@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        @a@�q�q�?             "@                        �a@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     "@	                        �a@)O���?             B@
                         �?�f7�z�?             =@            	          ����?���Q��?             4@                        �d@�n_Y�K�?	             *@                        0a@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     "@������������������������       �                     @�t�b�m0     h�h(h+K ��h-��R�(KMKK��h_�B0       �z@     �~@     �b@     �I@     �`@      4@     @X@       @     @W@      @     @V@      �?     �T@              @      �?              �?      @              @      @      �?      @      �?                      @      @              @      @       @      @       @                      @       @             �B@      (@      A@      @      ?@       @       @       @       @      �?       @                      �?              �?      7@              @      @      �?      @              @      �?               @              @      @       @      @              @       @      @      �?              �?      @      �?      �?      �?                      �?              @      �?              0@      ?@      (@      @              @      (@      @              �?      (@       @      (@      �?              �?      (@                      �?      @      9@      @      �?              �?      @                      8@     Pq@     �{@     �K@     Pw@       @     �`@      @     @]@      �?      �?              �?      �?              @      ]@      @     �\@             �U@      @      =@       @      &@       @      @      �?              �?      @              @      �?                       @      �?      2@              2@      �?               @      �?       @                      �?       @      1@       @      (@       @      @       @       @              �?       @      �?      �?              �?      �?              �?      �?                      @              @              @     �G@     �m@     �@@      N@       @      .@       @      �?              �?       @                      ,@      ?@     �F@      $@      ?@      $@      3@      @      2@      @      2@       @      2@               @       @      $@       @       @       @                       @               @       @              �?              @      �?      @                      �?              (@      5@      ,@      1@      ,@      @              *@      ,@      @              $@      ,@      $@      @      @              @      @       @      @              @       @       @       @                       @      @      �?              �?      @                      @      @              ,@     `f@      @      �?              �?      @              &@     @f@              >@      &@     �b@      @      @      @                      @       @     �a@       @     �^@       @      4@       @      @               @       @       @              �?       @      �?              �?       @                      0@      @     �Y@      @     �S@      @     �H@      @      G@      @      (@      �?      $@              @      �?      @              @      �?               @       @               @       @              �?      A@              7@      �?      &@      �?      �?      �?                      �?              $@       @      @       @                      @              =@              9@              3@     �k@     �P@      0@      8@      ,@      "@       @      "@       @       @              �?       @      �?       @                      �?              @      (@               @      .@      �?      .@               @      �?      @      �?                      @      �?             �i@     �E@     �g@      8@     �c@      .@      C@      "@      :@      "@      :@      @      @      @      �?      @      �?       @               @      �?                       @      @              6@       @      @       @      @                       @      0@                      @      (@             �]@      @      @       @      @                       @      ]@      @      ]@      @     @Q@             �G@      @      2@      @       @      @      @               @      @       @                      @      $@              =@                      �?      @@      "@      7@      "@      4@      @      *@      �?      *@                      �?      @       @       @       @      �?       @      �?      �?              �?      �?                      �?      �?              @              @      @      @       @      @                       @              @      "@              1@      3@      1@      (@       @      (@       @      @      @      @      @                      @      @                      @      "@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�\-hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�6         �       	          `ff�?��3����?A           ��@       C       
             �?*�����?2           �}@                           �?��a�n`�?e            `c@                           �J@���@M^�?             ?@                          `a@؇���X�?             5@                           �?�}�+r��?
             3@������������������������       �                     *@       	                   �n@r�q��?             @������������������������       �                     @
                          �d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                          �`@ףp=
�?             $@                          t@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @       *                    b@��� ��?Q             _@       )                    �? p�/��?6            @V@       "                   �[@ 	��p�?"             M@                           @O@�LQ�1	�?             7@                           �?      �?             0@              
             �?      �?              @������������������������       �                     @                          @_@z�G�z�?             @������������������������       �                     @              	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @        !       	          ����?����X�?             @������������������������       �                     @������������������������       �                      @#       $                    �O@��?^�k�?            �A@������������������������       �                     :@%       (                    `@�����H�?             "@&       '                    @P@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     ?@+       ,                    g@^������?            �A@������������������������       �        	             $@-       6                    �?�q�����?             9@.       /                    _@      �?              @������������������������       �                     @0       1                    @J@      �?             @������������������������       �                     �?2       3                   �b@�q�q�?             @������������������������       �                     �?4       5                   �c@      �?              @������������������������       �                     �?������������������������       �                     �?7       <                   �`@ҳ�wY;�?             1@8       9                    �?z�G�z�?             $@������������������������       �                     @:       ;                   �p@���Q��?             @������������������������       �                      @������������������������       �                     @=       >                   0a@և���X�?             @������������������������       �                     @?       B                   �a@      �?             @@       A       	            �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?D       O                   @E@�KM�]�?�            0t@E       N                    �?�n_Y�K�?             :@F       M       	            �?�\��N��?             3@G       J                    �?����X�?             ,@H       I                    �?      �?              @������������������������       �                     �?������������������������       �                     @K       L                     P@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @P       �                    �?�FVQ&�?�            �r@Q       h                    @L@~t�8��?�            `q@R       c       	             �?�h����?�             l@S       b                    �?`���˛?�            @k@T       a                    �?�x�V�?q             g@U       \                    �I@     ��?             @@V       W                    �?���7�?             6@������������������������       �                      @X       [                    l@P���Q�?
             4@Y       Z                   �e@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@]       ^                   �c@z�G�z�?             $@������������������������       �                     @_       `                    m@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        _             c@������������������������       �                    �@@d       g                   �_@r�q��?             @e       f                   Pn@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @i       j                   @Y@�����H�?!             K@������������������������       �                      @k       t                    �?$�q-�?              J@l       s       	          @33�?      �?              @m       n                    �L@      �?             @������������������������       �                     �?o       p                    �?�q�q�?             @������������������������       �                     �?q       r                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @u       v                    �?���7�?             F@������������������������       �                     9@w       x                    �?�KM�]�?             3@������������������������       �                     @y       z                   h@8�Z$���?
             *@������������������������       �                     @{       �                   �c@      �?              @|       }                   p@؇���X�?             @������������������������       �                     @~                            M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                   `_@D�n�3�?             3@������������������������       �                     @�       �                     N@և���X�?
             ,@�       �                   Pa@���!pc�?             &@������������������������       �                     �?�       �                    �?z�G�z�?             $@������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?NkL)���?           �{@�       �                    �?�q�q�?'            �P@�       �                    �?�p ��?            �D@�       �       	          033�?r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?��?^�k�?            �A@������������������������       �                     2@�       �                   `c@�IєX�?
             1@������������������������       �        	             0@������������������������       �                     �?�       �                    �?��H�}�?             9@�       �                   �r@�S����?             3@�       �                   �q@      �?             (@�       �                    �J@"pc�
�?
             &@�       �                   �V@      �?             @������������������������       �                     �?�       �                   �]@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �       
             �?\>ʆ4a�?�            `w@�       �                    �?     ��?�             t@�       �                    �R@�J��?�            �l@�       �                    �? (��?�            @l@�       �                   0j@�8��?n            �d@�       �                   �h@>a�����?#            �I@�       �                   Pe@���}<S�?              G@�       �                   @M@�X�<ݺ?             B@�       �       
             �?���}<S�?             7@�       �                   @\@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     4@������������������������       �                     *@�       �                    _@z�G�z�?             $@������������������������       �                     @�       �                   �f@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    @M@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                   0c@XB���?K             ]@�       �                    �J@����X�?H             \@�       �       	          `ff@ qP��B�?            �E@������������������������       �                    �A@�       �                    @J@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �        *            @Q@�       �       	          ����?      �?             @�       �                   �r@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �       	          ����?���#�İ?(            �M@�       �       
             �?�t����?             1@������������������������       �                      @������������������������       �        
             .@������������������������       �                     E@�       �                   �p@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                   P`@Z��:���?2            �V@�       �                    `@X�<ݚ�?             B@�       �                   �a@�g�y��?             ?@������������������������       �                     $@�       �                   �l@����X�?
             5@�       �                    �?ףp=
�?             $@������������������������       �                     @�       �                    �K@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    n@�eP*L��?             &@������������������������       �                     @�       �                   �c@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   b@�2����?            �K@������������������������       �                     C@�       �       	          ����?��.k���?             1@�       �       	          ����?؇���X�?             @�       �                   `^@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�z�G��?             $@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    �?��}*_��?             K@�       �                    @G@j���� �?             A@������������������������       �                     $@�       �                    �J@�q�q�?             8@������������������������       �                     @�       �                   �b@�\��N��?             3@�       �                   �b@���|���?             &@�       �       	          033�?      �?              @������������������������       �                     @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    e@      �?              @������������������������       �                     @������������������������       �                      @������������������������       �        	             4@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�       {@     P~@     @t@     @c@     �A@      ^@      3@      (@      2@      @      2@      �?      *@              @      �?      @              �?      �?      �?                      �?               @      �?      "@      �?      @              @      �?                      @      0@      [@      @     @U@      @      K@      @      4@      �?      .@      �?      @              @      �?      @              @      �?      �?              �?      �?                       @       @      @              @       @              �?      A@              :@      �?       @      �?       @      �?                       @              @              ?@      (@      7@              $@      (@      *@      @       @      @               @       @      �?              �?       @              �?      �?      �?      �?                      �?      @      &@       @       @              @       @      @       @                      @      @      @      @              �?      @      �?       @      �?                       @              �?     r@      A@      $@      0@      $@      "@      $@      @      @      �?              �?      @              @      @      @                      @              @              @     pq@      2@     �p@      $@     �k@      @     �j@      @     �f@      @      =@      @      5@      �?       @              3@      �?      @      �?      @                      �?      0@               @       @      @              �?       @               @      �?              c@             �@@              @      �?      �?      �?      �?                      �?      @              H@      @               @      H@      @      @       @       @       @      �?              �?       @              �?      �?      �?              �?      �?              @              E@       @      9@              1@       @      @              &@       @      @              @       @      @      �?      @               @      �?              �?       @                      �?      &@       @      @              @       @      @       @      �?               @       @               @       @              @             @[@     �t@      F@      6@     �A@      @      �?      @      �?                      @      A@      �?      2@              0@      �?      0@                      �?      "@      0@      @      0@      @      "@       @      "@       @       @              �?       @      �?              �?       @                      @      �?                      @      @             @P@     Ps@     �F@     0q@      0@     �j@      ,@     �j@      (@     `c@       @     �E@      @      E@       @      A@       @      5@       @      �?              �?       @                      4@              *@       @       @              @       @      @       @                      @      @      �?      @                      �?      @      \@      �?     �[@      �?      E@             �A@      �?      @              @      �?                     @Q@      @      �?      �?      �?              �?      �?               @               @     �L@       @      .@       @                      .@              E@       @      �?              �?       @              =@      O@      4@      0@      .@      0@              $@      .@      @      "@      �?      @              @      �?      @                      �?      @      @              @      @      �?              �?      @              @              "@      G@              C@      "@       @      @      �?      @      �?              �?      @              @              @      @      @       @      @                       @              @      4@      A@      4@      ,@      $@              $@      ,@              @      $@      "@      @      @      �?      @              @      �?      �?      �?                      �?      @              @       @      @                       @              4@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJI��$hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvMhwh(h+K ��h-��R�(KM��h~�B�8         �                    �?��e�B��?Q           ��@       ]                   �b@�G`N�"�?C           �@       >       
             �?|B���?           �y@                           �?@kT�3��?�            Pu@                          ``@^����?            �E@       	       	          ����?��.k���?
             1@                           a@z�G�z�?             $@������������������������       �                      @������������������������       �                      @
                           �?؇���X�?             @              	          ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                          p`@ȵHPS!�?             :@              	             �?d}h���?
             ,@                           ^@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     (@       ;                    �R@@c`�}y�?�            �r@                          �U@�;��m��?�            `r@������������������������       �                      @       (                    @G@�V����?�            @r@                           �?�q��/��?            �H@������������������������       �                     &@       '       	          033@�S����?             C@       &       	          ����?�����H�?             B@       #                   Pg@�㙢�c�?             7@       "                    �D@�q�q�?             "@        !                    �C@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @$       %                    �?@4և���?             ,@������������������������       �                     *@������������������������       �                     �?������������������������       �        	             *@������������������������       �                      @)       .       	          ����? ��u좤?�            `n@*       +       	          ����?��<D�m�?             �H@������������������������       �                     F@,       -                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @/       2                   �Q@�a�O�?{            @h@0       1                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?3       :                   �N@�f]/U�?y            �g@4       5                   �]@ qP��B�?            �E@������������������������       �                     4@6       9                   @^@�nkK�?             7@7       8                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     3@������������������������       �        ^            �b@<       =                   �p@      �?             @������������������������       �                      @������������������������       �                      @?       L                    �?��.k���?0             Q@@       E                    �?�I�w�"�?             C@A       D                    P@ �q�q�?             8@B       C       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     6@F       K                   `@և���X�?             ,@G       J                     K@z�G�z�?             $@H       I       	          ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @M       R       	             �?�������?             >@N       Q                   e@X�<ݚ�?             "@O       P                   0a@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @S       T                   �_@؇���X�?             5@������������������������       �                     &@U       \                   `W@�z�G��?             $@V       W                    �?      �?             @������������������������       �                      @X       [                    �?      �?             @Y       Z                   `b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @^       m                    k@�"���r�?;            �X@_       l                    �?��hJ,�?             A@`       c                    �E@���N8�?             5@a       b       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @d       e                   Pc@r�q��?	             2@������������������������       �                     �?f       g                   @[@�t����?             1@������������������������       �                     �?h       i                   `@      �?             0@������������������������       �                     $@j       k                   �d@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             *@n              
             �?�G\�c�?&            @P@o       t                     M@�5��?             ;@p       q                   �r@�C��2(�?             &@������������������������       �                     @r       s                    �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @u       v       
             �?      �?	             0@������������������������       �                     �?w       ~                    �?�q�q�?             .@x       }       	             @r�q��?             (@y       |                   �r@�C��2(�?             &@z       {                   �q@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   Pd@p9W��S�?             C@�       �                   �_@և���X�?             5@�       �                    �?"pc�
�?             &@������������������������       �                      @������������������������       �                     "@������������������������       �                     $@�       �                     N@�t����?             1@�       �                   `a@      �?
             0@������������������������       �                     &@�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   �q@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �       
             �?�������?           �y@�       �                    @F@`n��k��?c            `a@�       �                   (p@ףp=
�?             4@�       �                    �?�}�+r��?             3@������������������������       �                     0@�       �                   �l@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �       
             �?<����l�?T            �]@�       �                   `a@�n_Y�K�?             *@�       �                    �?����X�?             @������������������������       �                     �?�       �                    b@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	          ����?r�0p�?H            �Z@�       �                    �?�>����?             ;@�       �                   �h@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @M@ �q�q�?             8@�       �                    �K@�C��2(�?	             &@������������������������       �                     "@�       �                   0a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             *@�       �                   �b@v�_���?3            �S@�       �                   p`@@�0�!��?"            �I@�       �                    k@j���� �?             1@�       �                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                   �^@���Q��?	             $@�       �       	          033�?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @N@r�q��?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�IєX�?             A@������������������������       �                     �?�       �                   �`@Pa�	�?            �@@������������������������       �                     7@�       �                   �a@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�       �                   (p@X�Cc�?             <@�       �                    �K@r�q��?             2@�       �                    �?�q�q�?             "@������������������������       �                     @�       �                   �K@      �?             @������������������������       �                      @�       �                   �c@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@�       �       	          ����?�z�G��?             $@�       �                   �c@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�                         @g@��j���?�            �p@�       �                    @L@�)2e��?�            �p@�       �                    @�k~X��?�             k@�       �       	          ���@���9�,�?|             i@�       �                   c@@��d�`�?{             i@�       �                   @[@ ��N8�?7             U@�       �                    �E@؇���X�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        3            @S@������������������������       �        D             ]@������������������������       �                     �?�       �                    �?��S�ۿ?             .@������������������������       �                     ,@������������������������       �                     �?�             	          `ff�?�c�����?'            �J@�       �                    c@r�q��?$             H@�       �                    @M@��-�=��?            �C@�       �                    �?�θ�?	             *@�       �                    �?և���X�?             @������������������������       �                     �?�       �                   �a@�q�q�?             @������������������������       �                     @�       �                   0b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          ����? ��WV�?             :@�       �                    �O@�8��8��?	             (@������������������������       �                      @�       �                   �r@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             ,@�                            R@X�<ݚ�?             "@�       �                   �k@����X�?             @������������������������       �                      @�       �       	          ����?���Q��?             @�       �                   �`@�q�q�?             @������������������������       �                     �?�       �                   �m@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KMKK��h_�B0       �y@     �@     �Z@      y@     �O@     �u@      ;@     �s@      (@      ?@      "@       @       @       @       @                       @      �?      @      �?      �?              �?      �?                      @      @      7@      @      &@      @      @              @      @                       @              (@      .@     �q@      *@     �q@       @              &@     �q@      @     �E@              &@      @      @@      @      @@      @      3@      @      @      @       @               @      @                      @      �?      *@              *@      �?                      *@       @              @     �m@      @      G@              F@      @       @      @                       @       @      h@      �?       @               @      �?              �?     �g@      �?      E@              4@      �?      6@      �?      @              @      �?                      3@             �b@       @       @               @       @              B@      @@      =@      "@      7@      �?      �?      �?      �?                      �?      6@              @       @       @       @       @      �?              �?       @                      @      @              @      7@      @      @      @       @               @      @                      @      @      2@              &@      @      @      @      @       @              �?      @      �?      �?              �?      �?                       @              @     �E@      L@      @      =@      @      0@       @      �?              �?       @              @      .@      �?               @      .@      �?              �?      .@              $@      �?      @              @      �?                      *@      C@      ;@      &@      0@      �?      $@              @      �?      @      �?                      @      $@      @              �?      $@      @      $@       @      $@      �?      @      �?      @                      �?      @                      �?              @      ;@      &@      (@      "@       @      "@       @                      "@      $@              .@       @      .@      �?      &@              @      �?       @               @      �?       @                      �?              �?     @s@     �Y@     �K@      U@      2@       @      2@      �?      0@               @      �?       @                      �?              �?     �B@     �T@       @      @       @      @      �?              �?      @              @      �?              @              =@     @S@       @      9@      �?       @      �?                       @      �?      7@      �?      $@              "@      �?      �?      �?                      �?              *@      ;@      J@      "@      E@      @      $@      �?      @      �?                      @      @      @      �?      @               @      �?      �?      �?                      �?      @      �?      @              �?      �?              �?      �?               @      @@      �?              �?      @@              7@      �?      "@      �?                      "@      2@      $@      .@      @      @      @      @              @      @               @      @      �?              �?      @              "@              @      @      @       @      @                       @              @     �o@      2@     �o@      0@     �j@      @     �h@       @     �h@      �?     �T@      �?      @      �?      @              �?      �?      �?                      �?     @S@              ]@                      �?      ,@      �?      ,@                      �?      D@      *@      D@       @     �A@      @      $@      @      @      @              �?      @       @      @              �?       @               @      �?              @              9@      �?      &@      �?       @              @      �?      @                      �?      ,@              @      @      @       @       @              @       @      �?       @              �?      �?      �?              �?      �?               @                       @              @               @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���;hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM	hwh(h+K ��h-��R�(KM	��h~�B�9         �       
             �?�5�C��?@           ��@       s                   �b@�N��R��?G           ��@                           �?L��n��?           �{@                           �?      �?"             K@                           �?�n_Y�K�?            �C@              	             �?     ��?             @@                           �B@l��[B��?             =@������������������������       �                     @	                           �?      �?             8@
                          �`@և���X�?             5@������������������������       �                      @                          pb@�	j*D�?             *@������������������������       �                     @                            L@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @                           �?z�G�z�?
             .@������������������������       �                      @                          Hp@�θ�?	             *@������������������������       �                     "@                          �`@      �?             @                          @_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @       >                    �?���2"��?�             x@       #       	          ����?��j���??            �[@                            �K@����?�?            �F@������������������������       �                     =@!       "                   �X@      �?             0@������������������������       �                     �?������������������������       �                     .@$       3                    �?r٣����?'            �P@%       &                     G@���|���?            �@@������������������������       �                     @'       (                   �^@�c�Α�?             =@������������������������       �                     @)       .                   �k@���|���?             6@*       +                    �K@�eP*L��?             &@������������������������       �                     @,       -                   �b@؇���X�?             @������������������������       �                     @������������������������       �                     �?/       0                   @_@"pc�
�?             &@������������������������       �                     @1       2                    �?����X�?             @������������������������       �                     @������������������������       �                      @4       9                    �?<���D�?            �@@5       6       	          ����?�q�q�?             @������������������������       �                     �?7       8                   `c@      �?              @������������������������       �                     �?������������������������       �                     �?:       =                   `R@��S�ۿ?             >@;       <                    Q@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ;@?       J                   `_@���!���?�            0q@@       I                    \@X;��?i            @f@A       F       	             �?(a��䛼?:            @Y@B       C       	          ����?�r����?             >@������������������������       �                     9@D       E                   �Y@z�G�z�?             @������������������������       �                     �?������������������������       �                     @G       H                    `R@�J�T�?(            �Q@������������������������       �        '            @Q@������������������������       �                      @������������������������       �        /            @S@K       j       	          `ff�?��l��?B            @X@L       i                   �n@D>�Q�?&             J@M       `                    �?���"͏�?            �B@N       S                    �D@r�q��?             >@O       P       	             �?և���X�?             @������������������������       �                     @Q       R                   g@      �?             @������������������������       �                     @������������������������       �                     �?T       Y                   �_@���}<S�?             7@U       X                    �?      �?             @V       W                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @Z       [                   `a@�}�+r��?             3@������������������������       �                     (@\       _                    b@؇���X�?             @]       ^                    ^@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @a       b       	             �?և���X�?             @������������������������       �                     �?c       d                   f@�q�q�?             @������������������������       �                     �?e       f                    �?z�G�z�?             @������������������������       �                     �?g       h                   Pb@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     .@k       r                   `j@`Ӹ����?            �F@l       o                   �i@؇���X�?
             ,@m       n                   �U@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@p       q                   �^@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ?@t       �                    �M@z�J��?;            �W@u       z                    �?�e����?/            �S@v       y                   q@��2(&�?             6@w       x       	          ���@P���Q�?             4@������������������������       �                     3@������������������������       �                     �?������������������������       �                      @{       �                    �?~h����?"             L@|       �                   �r@     ��?             0@}       ~                   �k@�r����?
             .@������������������������       �                      @       �                   `q@����X�?             @�       �                    �F@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    @���Q��?             D@�       �       	          ����?r֛w���?             ?@�       �                    �?և���X�?             @�       �                   �_@      �?             @������������������������       �                      @�       �                    �E@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                     G@r�q��?             8@������������������������       �                     *@�       �                   �h@���|���?             &@������������������������       �                      @�       �                   @d@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    �?�����H�?             "@�       �                   @b@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?�       �                   xu@      �?             0@�       �       	          `ff@@4և���?
             ,@������������������������       �                     &@�       �       
             �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                   pc@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?     N�?�             x@�       �                    @L@�MI8d�?�            �t@�       �                   @E@���>�?�            �n@�       �                   �\@������?
             .@������������������������       �                      @�       �                   �c@8�Z$���?             *@�       �                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�       �                    �? :��?�            �l@�       �                     I@"pc�
�?            �@@�       �                   0f@�q�q�?
             .@������������������������       �                     @������������������������       �                     $@�       �                    g@�X�<ݺ?             2@������������������������       �                     1@������������������������       �                     �?�       �                    �?`�LVXz�?�            �h@�       �                    �? h'M#�?{            �f@�       �                    @I@�7��?            �C@������������������������       �                     ;@�       �                   �d@r�q��?             (@�       �                   Pm@�C��2(�?             &@�       �                    ]@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?������������������������       �        c             b@������������������������       �        	             .@�       �       	          `ff�?|�|k6��?5            �U@�       �                    @�q�q�?.            �S@�       �                   �b@4�	~���?)            @Q@�       �                   @_@:�&���?            �C@�       �                   @Z@��
ц��?             *@������������������������       �                     @�       �                    �?؇���X�?             @�       �                    ^@      �?             @�       �                    �P@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                   �_@ ��WV�?             :@�       �                   �^@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@�       �                   �q@      �?             >@�       �                    @M@�	j*D�?	             *@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�����H�?             "@������������������������       �                     @�       �                    �?      �?             @�       �                   �c@�q�q�?             @������������������������       �                     �?�       �                   �i@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �       	          ����?ҳ�wY;�?
             1@�       �                    �?d}h���?             ,@�       �                    �?�C��2(�?             &@�       �                    s@      �?              @�       �                   �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                   @`@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                     "@�                         Pd@��.k���?             �I@�       �                   Pj@�zv�X�?             F@�       �                    `@���y4F�?             3@������������������������       �                     @�       �                   �`@�q�q�?             (@�       �       	          033�?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�                          �L@�q�����?             9@�                           �H@r�q��?             (@�       �                   0a@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     "@                        �_@�θ�?	             *@                         b@      �?              @                         [@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM	KK��h_�B�       �y@     �@     @[@     �z@     �N@     �w@      ;@      ;@      .@      8@      .@      1@      .@      ,@              @      .@      "@      (@      "@       @              @      "@              @      @      @      @                      @      @                      @              @      (@      @       @              $@      @      "@              �?      @      �?      �?              �?      �?                       @      A@      v@      1@     �W@      �?      F@              =@      �?      .@      �?                      .@      0@      I@      (@      5@      @               @      5@              @       @      ,@      @      @              @      @      �?      @                      �?       @      "@              @       @      @              @       @              @      =@       @      �?      �?              �?      �?      �?                      �?       @      <@       @      �?              �?       @                      ;@      1@      p@      @     �e@      @     �W@      @      :@              9@      @      �?              �?      @               @     @Q@             @Q@       @                     @S@      &@     �U@      "@     �E@      "@      <@      @      9@      @      @              @      @      �?      @                      �?       @      5@      �?      @      �?      �?      �?                      �?               @      �?      2@              (@      �?      @      �?      @      �?                      @               @      @      @              �?      @       @              �?      @      �?      �?              @      �?      @                      �?              .@       @     �E@       @      (@      �?      &@      �?                      &@      �?      �?      �?                      �?              ?@      H@      G@      G@      @@      3@      @      3@      �?      3@                      �?               @      ;@      =@      @      *@       @      *@               @       @      @       @      �?              �?       @                      @      �?              8@      0@      7@       @      @      @      @      �?       @              �?      �?      �?                      �?              @      4@      @      *@              @      @               @      @       @      @                       @      �?       @      �?      @              @      �?                      �?       @      ,@      �?      *@              &@      �?       @               @      �?              �?      �?              �?      �?             �r@     @T@     pq@      K@     `l@      3@      @      &@       @               @      &@       @      @              @       @                       @     �k@       @      ;@      @      $@      @              @      $@              1@      �?      1@                      �?     �h@       @     �f@       @     �B@       @      ;@              $@       @      $@      �?      @      �?              �?      @              @                      �?      b@              .@              J@     �A@      J@      :@     �G@      6@      @@      @      @      @      @              �?      @      �?      @      �?      �?              �?      �?                       @              @      9@      �?      @      �?      @                      �?      2@              .@      .@      "@      @      �?      @              @      �?               @      �?      @              @      �?       @      �?      �?              �?      �?              �?      �?              �?              @      &@      @      &@      �?      $@      �?      @      �?      @              @      �?                      @              @       @      �?       @                      �?      @              @      @              @      @                      "@      8@      ;@      1@      ;@      @      .@              @      @       @      @      @              @      @                      @      *@      (@      $@       @      �?       @      �?                       @      "@              @      $@      @      @      @      �?              �?      @                      @              @      @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�n�KhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM'hwh(h+K ��h-��R�(KM'��h~�B�@         �                   �`@���3L�?7           ��@                           �?*)ώ-��?           �z@                           �?�[�IJ�?!            �G@                          �R@�E��ӭ�?             B@������������������������       �                      @                          �s@������?             A@                           b@؇���X�?             <@       	                   Xp@���}<S�?             7@������������������������       �                     0@
                           �O@����X�?             @                          @[@���Q��?             @                           �?�q�q�?             @                          `X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @                           �O@���Q��?             @������������������������       �                     @������������������������       �                      @              	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     @              	             �?�C��2(�?             &@                           �O@      �?             @              
             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @        U                    �?�/z���?�            �w@!       P       	          ����?~�u���?]            �a@"       1                    @K@r�q��?C             X@#       $                    @A@�q�q�?             E@������������������������       �                      @%       .                    �?�z�G��?             D@&       -       
             �?      �?             6@'       ,                    �?�8��8��?	             (@(       +                    �I@      �?             @)       *       	             �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     $@/       0                    �?�X�<ݺ?             2@������������������������       �                     �?������������������������       �                     1@2       G       
             �?�E��ӭ�?%             K@3       F                   �v@�KM�]�?             C@4       C                    @�L���?            �B@5       6                   �W@�FVQ&�?            �@@������������������������       �                     "@7       <                    @L@�8��8��?             8@8       ;                    �?z�G�z�?             @9       :                   �X@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @=       B                    �?�}�+r��?             3@>       ?                    �O@ףp=
�?             $@������������������������       �                      @@       A                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@D       E                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?H       K                    �?     ��?             0@I       J                   �\@�q�q�?             @������������������������       �                      @������������������������       �                     @L       O                    �?ףp=
�?             $@M       N                   �n@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @Q       R                    �Q@=QcG��?            �G@������������������������       �                     D@S       T                    �?և���X�?             @������������������������       �                     @������������������������       �                     @V       }                    �?p�U�ʻ�?�            �m@W       f       	          hff�?(a��䛼?x            @i@X       c                   (p@     ��?             @@Y       b                    �?@4և���?             <@Z       [                    �M@$�q-�?             :@������������������������       �                     (@\       a                    �?؇���X�?             ,@]       ^                    �?�<ݚ�?             "@������������������������       �                     @_       `       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @d       e                    b@      �?             @������������������������       �                     @������������������������       �                     �?g       h                    @J@h�|�6�?c            @e@������������������������       �                    �H@i       n                   �h@��a��?H            @^@j       k                    c@@��8��?             H@������������������������       �                     C@l       m                   @`@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?o       x                   ``@�F��O�?,            @R@p       s       	          ����?z�G�z�?             9@q       r                    �?      �?             @������������������������       �                     @������������������������       �                     �?t       u       	          033@�����?             5@������������������������       �                     2@v       w                    �J@�q�q�?             @������������������������       �                      @������������������������       �                     �?y       |       
             �?@��8��?             H@z       {                   �c@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     F@~                           Y@��G���?            �B@������������������������       �                     @�       �                    @�t����?             A@�       �       	          ����?     ��?             @@�       �                   p`@      �?             (@�       �                    �?      �?             @�       �                    `P@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     4@�       �                   �j@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       	          ����?�%���h�?+           �~@�       �                   @E@ ��3��?�            pr@�       �                   �Y@@4և���?
             ,@������������������������       �                     �?������������������������       �        	             *@�       �                   pq@@�"[R&�?�            �q@�       �                    �?v`N����?�            �k@�       �       	          ����?t�U����?{             i@�       �       
             �?�׾���?w             h@�       �                   0e@J�8���?             =@�       �       	          ����?��<b���?             7@�       �                    �?և���X�?             @������������������������       �                     @������������������������       �                     @�       �                    �?      �?             0@�       �                    �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?$�q-�?             *@������������������������       �                      @�       �                   pn@z�G�z�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   n@r�q��?             @������������������������       �                     @�       �                   �n@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @L@0��P�?e            �d@�       �                    �?�lm�9�?X            �a@�       �                   �i@     ��?             @@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @D@ 	��p�?             =@�       �                    a@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �l@ 7���B�?
             ;@������������������������       �                     1@�       �                    �?ףp=
�?             $@������������������������       �                     �?�       �                   `m@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                   @[@��wڝ�?I            @[@�       �                    m@�C��2(�?             &@������������������������       �                      @�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        B            �X@�       �                    �N@��+7��?             7@�       �                    �?��
ц��?             *@������������������������       �                     @�       �                    �L@      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     $@�       �                    �H@      �?              @������������������������       �                     @������������������������       �                     @�       �                   �b@      �?             6@�       �                   �`@"pc�
�?             &@������������������������       �                     �?�       �                    �J@ףp=
�?             $@�       �       
             �?      �?             @������������������������       �                     �?�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?"pc�
�?	             &@������������������������       �                     @�       �                    �?���Q��?             @������������������������       �                      @������������������������       �                     @�       �       
             �?J�8���?#             M@�       �                    @O@�IєX�?
             1@������������������������       �        	             0@������������������������       �                     �?�       �                   Pe@������?            �D@�       �                    �?@-�_ .�?            �B@�       �                    �M@8�Z$���?             *@������������������������       �                     $@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     8@�       �                    �?      �?             @�       �                   f@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�             	          ���@�E���?r            @h@�                          �?z�J��?U            �a@�       �                   `Y@rp��P��?1            �T@������������������������       �                     @�                         xr@�G�z.�?/             T@�       �                    �?��M���?(             Q@�       �       	          033�?�}�+r��?
             3@�       �                    �L@      �?              @�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�       �                    @F@f�Sc��?            �H@������������������������       �                     $@�       �                     I@��
ц��?            �C@������������������������       �                      @                         Hq@�4�����?             ?@                        �b@�<ݚ�?             ;@      	      	          ����?"pc�
�?             6@            	             �?և���X�?             @                         �?�q�q�?             @������������������������       �                     �?                          @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?
                         �?��S�ۿ?	             .@������������������������       �                     �?������������������������       �                     ,@            
             �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     (@                        �l@\-��p�?$             M@                        e@������?             >@                        �k@d}h���?             <@                        Pg@�8��8��?             8@                         �?z�G�z�?             $@                         �G@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     ,@������������������������       �                     @������������������������       �                      @������������������������       �                     <@      $                   �F@ �h�7W�?            �J@       !      	          033@"pc�
�?             &@������������������������       �                     @"      #                  pk@���Q��?             @������������������������       �                      @������������������������       �                     @%      &                  �e@�Ń��̧?             E@������������������������       �                    �D@������������������������       �                     �?�t�b��0     h�h(h+K ��h-��R�(KM'KK��h_�Bp       px@     x�@      W@     u@      ;@      4@      :@      $@               @      :@       @      8@      @      5@       @      0@              @       @      @       @      �?       @      �?      �?              �?      �?                      �?       @               @              @       @      @                       @       @      @       @                      @      �?      $@      �?      @      �?      �?              �?      �?                       @              @     @P@     �s@      G@     @X@     �E@     �J@      <@      ,@               @      <@      (@      &@      &@      �?      &@      �?      @      �?      �?              �?      �?                       @               @      $@              1@      �?              �?      1@              .@     �C@      @      A@      @      A@       @      ?@              "@       @      6@      �?      @      �?      �?      �?                      �?              @      �?      2@      �?      "@               @      �?      �?              �?      �?                      "@      �?      @              @      �?              �?              &@      @       @      @       @                      @      "@      �?      @      �?      @                      �?      @              @      F@              D@      @      @              @      @              3@     �k@      (@     �g@      @      ;@       @      :@       @      8@              (@       @      (@       @      @              @       @      �?              �?       @                      @               @      @      �?      @                      �?      @     `d@             �H@      @     �\@      �?     �G@              C@      �?      "@              "@      �?              @     �P@      @      4@      @      �?      @                      �?       @      3@              2@       @      �?       @                      �?      �?     �G@      �?      @              @      �?                      F@      @      >@      @              @      >@      @      =@      @      "@      @      @      @       @      @                       @              �?              @              4@      �?      �?      �?                      �?     �r@     �g@     `l@      Q@      �?      *@      �?                      *@     @l@     �K@     �g@     �A@      f@      8@     �e@      4@      3@      $@      2@      @      @      @              @      @              ,@       @       @      �?              �?       @              (@      �?       @              @      �?      �?      �?              �?      �?              @              �?      @              @      �?       @      �?                       @     @c@      $@      a@      @      =@      @       @      �?              �?       @              ;@       @      �?      �?      �?                      �?      :@      �?      1@              "@      �?      �?               @      �?              �?       @              [@      �?      $@      �?       @               @      �?       @                      �?     �X@              1@      @      @      @              @      @      �?       @      �?              �?       @              @              $@              @      @      @                      @      &@      &@       @      "@      �?              �?      "@      �?      @              �?      �?       @               @      �?                      @      "@       @      @              @       @               @      @              C@      4@      �?      0@              0@      �?             �B@      @     �A@       @      &@       @      $@              �?       @               @      �?              8@               @       @      �?       @               @      �?              �?              R@     �^@     @Q@      R@     �N@      6@              @     �N@      3@     �H@      3@      2@      �?      @      �?      �?      �?      �?                      �?      @              &@              ?@      2@      $@              5@      2@               @      5@      $@      5@      @      2@      @      @      @      @       @              �?      @      �?      @                      �?              �?      ,@      �?              �?      ,@              @       @               @      @                      @      (@               @      I@       @      6@      @      6@       @      6@       @       @       @      �?              �?       @                      @              ,@      @               @                      <@      @      I@       @      "@              @       @      @       @                      @      �?     �D@             �D@      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���-hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK�h~�B�4         4                    `@�$�����?I           ��@                           �?����M�?l            �e@              
             �?��sK�z�?N            �^@                           @K@���!pc�?             &@                            H@�q�q�?             @������������������������       �                     �?������������������������       �                      @       	                   @\@      �?              @������������������������       �                     @
                           �?      �?              @������������������������       �                     �?������������������������       �                     �?              	          033�?h�����?G             \@              
             �?�}��L�?0            �R@������������������������       �        %             K@                           @I@���N8�?             5@������������������������       �                     $@                           �J@�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@                           �?�L���?            �B@                           �?(;L]n�?             >@              
             �?�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     2@                           �N@����X�?             @                          �a@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @        3                    �? �o_��?             I@!       0       
             �?��S���?             >@"       '                    �?�LQ�1	�?             7@#       &                    �?z�G�z�?	             .@$       %                   �\@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@(       -                    �?      �?              @)       *       	          `ff�?      �?             @������������������������       �                     �?+       ,                     @�q�q�?             @������������������������       �                      @������������������������       �                     �?.       /                   �b@      �?             @������������������������       �                     �?������������������������       �                     @1       2                    `Q@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �        
             4@5       z                   a@Һ9���?�           H�@6       s       
             �?;��1��?�             t@7       b                   Xs@���ʂ��?�            �n@8       C                    �?LܤK���?�            �j@9       :                    _@�eP*L��?             6@������������������������       �                     @;       B                    `P@      �?             0@<       =                   @]@�θ�?
             *@������������������������       �                     @>       A                   �`@և���X�?             @?       @                   �_@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @D       I                     E@p�q��?t             h@E       F                    @D@�z�G��?             $@������������������������       �                     @G       H                    �?      �?             @������������������������       �                     @������������������������       �                     �?J       U                   �[@�ȉo(��?m            �f@K       N                   @\@���;QU�?(            @R@L       M                     O@�q�q�?             @������������������������       �                     @������������������������       �                      @O       P                   @a@�����?$            �P@������������������������       �                     @@Q       R                   `[@�#-���?            �A@������������������������       �                     =@S       T                    �L@      �?             @������������������������       �                     @������������������������       �                     @V       a                    �?бK/eh�?E            @[@W       `                   �r@ �Cc}�?             <@X       Y                     O@�>����?             ;@������������������������       �                     2@Z       _                     P@�<ݚ�?             "@[       \                   0k@���Q��?             @������������������������       �                      @]       ^       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �        4            @T@c       d                    T@���!pc�?            �@@������������������������       �                      @e       r                   �e@��a�n`�?             ?@f       g                    �?д>��C�?             =@������������������������       �                      @h       o                   ``@���N8�?             5@i       n                    �?և���X�?             @j       k                    ]@z�G�z�?             @������������������������       �                     �?l       m                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @p       q       
             �?؇���X�?
             ,@������������������������       �                      @������������������������       �        	             (@������������������������       �                      @t       y       	             �?`2U0*��?/            �R@u       v                    �? �й���?-            @R@������������������������       �        '             P@w       x                   �b@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                      @{       �       
             �?p�v>��?           pz@|       �                   �o@
j*D>�?j            �c@}       �                    �?4���C�??            �X@~              
             �?��R[s�?            �A@������������������������       �                     $@�       �                     F@��H�}�?             9@������������������������       �                     @�       �                   �b@�\��N��?             3@�       �                    �M@X�Cc�?             ,@�       �       	          ����?      �?	             (@�       �                   �_@�q�q�?             "@������������������������       �                      @�       �       	             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   `a@      �?)             P@�       �                    @L@�iʫ{�?!            �J@�       �                    �?$�q-�?            �C@�       �                    �?�g�y��?             ?@�       �       
             �?�C��2(�?             &@�       �                   �\@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �                     4@�       �                   0d@      �?              @������������������������       �                      @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    �?և���X�?             ,@�       �       	          033@�q�q�?             "@�       �       	          ����?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �       	          033�?���|���?             &@�       �                   pk@؇���X�?             @������������������������       �                     @�       �                    �L@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?�S����?+            �L@�       �                    �?��X��?             <@�       �                   �b@      �?             8@�       �       	          ����?�G�z��?             4@�       �       	          ����?X�Cc�?             ,@�       �                    �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     =@�       �                    �?4�<����?�            �p@�       �                    �?�E��
��?%             J@�       �                   �j@�f7�z�?             =@������������������������       �                     @�       �                   ``@
;&����?             7@�       �                   �c@      �?
             0@������������������������       �                     @�       �                    �?���Q��?             $@�       �                   �d@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �                    �J@      �?             @������������������������       �                      @������������������������       �                      @�       �                    �?؇���X�?             @�       �                   �b@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                     L@�㙢�c�?             7@������������������������       �                     *@�       �                   `c@���Q��?             $@�       �                   �d@      �?              @�       �                    �?z�G�z�?             @������������������������       �                      @�       �                    w@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                   `]@Du9iH��?�            �j@�       �                   �l@z�G�z�?            �F@������������������������       �                     4@�       �                   �l@��H�}�?             9@������������������������       �                     @�       �                   @[@�S����?             3@�       �                   @c@�q�q�?             @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    @N@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?�       �                    �?@�)�n�?m            @e@�       �                     I@b�h�d.�?            �A@������������������������       �                     6@�       �                    @J@��
ц��?
             *@������������������������       �                     @�       �       	             �?�z�G��?             $@�       �                   pc@      �?              @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �        U            �`@�t�bh�h(h+K ��h-��R�(KK�KK��h_�B       `z@      @      5@      c@      @      ]@      @       @       @      �?              �?       @              �?      @              @      �?      �?      �?                      �?      @      [@      �?     �R@              K@      �?      4@              $@      �?      $@      �?                      $@      @      A@      �?      =@      �?      &@              &@      �?                      2@       @      @       @      �?       @                      �?              @      ,@      B@      ,@      0@       @      .@      @      (@      @       @      @                       @              $@      @      @       @       @              �?       @      �?       @                      �?      @      �?              �?      @              @      �?      @                      �?              4@     y@     �u@      Z@     @k@      @@     �j@      7@     �g@      (@      $@      @              @      $@      @      $@              @      @      @      @      �?      @                      �?              @      @              &@     �f@      @      @              @      @      �?      @                      �?       @     �e@      @      Q@       @      @              @       @              @      P@              @@      @      @@              =@      @      @      @                      @      @     �Z@      @      9@       @      9@              2@       @      @       @      @               @       @      �?              �?       @                      @      �?                     @T@      "@      8@       @              @      8@      @      8@               @      @      0@      @      @      �?      @              �?      �?      @      �?                      @       @               @      (@       @                      (@       @              R@      @      R@      �?      P@               @      �?       @                      �?               @     �r@     �_@     �P@     �V@     �L@      E@      "@      :@              $@      "@      0@              @      "@      $@      "@      @      "@      @      @      @               @      @      �?      @                      �?      @                       @              @      H@      0@      F@      "@      B@      @      >@      �?      $@      �?      �?      �?              �?      �?              "@              4@              @       @       @              @       @               @      @               @      @      @      @      @       @               @      @                      @      @              @      @      �?      @              @      �?      �?              �?      �?              @      �?      @                      �?      "@      H@      "@      3@      "@      .@      "@      &@      "@      @      �?      @      �?                      @       @                      @              @              @              =@     �l@      B@      ?@      5@      (@      1@              @      (@      &@      @      $@              @      @      @      @       @      @                       @       @       @       @                       @      @      �?       @      �?       @                      �?      @              3@      @      *@              @      @      @      @      �?      @               @      �?       @               @      �?              @               @              i@      .@      B@      "@      4@              0@      "@              @      0@      @      @       @      �?       @      �?                       @      @              (@      �?      (@                      �?     �d@      @      =@      @      6@              @      @              @      @      @      @      �?      @               @      �?              �?       @                       @     �`@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ���hG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�7         �       
             �?�HK��x�?O           ��@       �                    �R@w�)_��?L           �@       r                   �b@b<g���?K           �@              	          ����?��,��?           �{@������������������������       �        7            @X@              	          ����?d	��g��?�            �u@       
                   @b@և���X�?             ,@       	                    @I@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @                           @I@z�G�z�?             @������������������������       �                     �?������������������������       �                     @       1                    �?H�q�R��?�            �t@                           �?V������?/            �R@                          �`@�q�q�?             5@                          `X@؇���X�?
             ,@������������������������       �                     �?                           @L@$�q-�?	             *@              	             �?r�q��?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @                           �?����X�?             @������������������������       �                     @������������������������       �                      @       0                   pe@f1r��g�?"            �J@       #       	             �?�t����?!            �I@               
             �?���Q��?             @������������������������       �                      @!       "       	          033�?�q�q�?             @������������������������       �                     �?������������������������       �                      @$       /                    �?���.�6�?             G@%       &                    �?ܷ��?��?             =@������������������������       �                     &@'       .       	          `ff�?r�q��?             2@(       )       
             �?�q�q�?             "@������������������������       �                     �?*       +                    �G@      �?              @������������������������       �                      @,       -                   `@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     "@������������������������       �        
             1@������������������������       �                      @2       C                    �?����?�            Pp@3       @                   @b@���!pc�?             6@4       5                   @_@      �?             0@������������������������       �                     @6       9       	          ����?z�G�z�?	             $@7       8                    @O@      �?              @������������������������       �                     �?������������������������       �                     �?:       ?                   ``@      �?              @;       >                    �?�q�q�?             @<       =                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @A       B                   `^@�q�q�?             @������������������������       �                      @������������������������       �                     @D       Y       	          ����?��'���?�            �m@E       J       	          `ff�?��v����?)            �P@F       G                   �j@���7�?             6@������������������������       �        
             2@H       I                   �`@      �?             @������������������������       �                     @������������������������       �                     �?K       N                   �[@:	��ʵ�?            �F@L       M                    `@�q�q�?             @������������������������       �                     �?������������������������       �                      @O       V                    �?؇���X�?             E@P       U                   �X@Pa�	�?            �@@Q       R                    �K@�����H�?             "@������������������������       �                     @S       T                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     8@W       X                   �l@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @Z       g                   �_@��+��<�?v            �e@[       d                   �c@�r�MȢ?M            �Z@\       c                   @_@��K2��?D            �W@]       ^                   po@���7�?             6@������������������������       �                     .@_       b                    �J@؇���X�?             @`       a                   @]@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        3             R@e       f                     R@$�q-�?	             *@������������������������       �                     (@������������������������       �                     �?h       q                    �J@����?)            @P@i       l                    `@"pc�
�?             6@j       k                   Ph@���Q��?             @������������������������       �                      @������������������������       �                     @m       p                    �?�t����?	             1@n       o                   �U@      �?             0@������������������������       �                     �?������������������������       �                     .@������������������������       �                     �?������������������������       �                    �E@s       �                    �?$/����?0            @P@t       �       	          ���@     ��?             @@u       v                    @L@V�a�� �?             =@������������������������       �                     .@w       x                    �L@և���X�?             ,@������������������������       �                     @y       �                    �?���!pc�?             &@z       }                    �?z�G�z�?             $@{       |                   pc@      �?              @������������������������       �                     �?������������������������       �                     �?~                          �c@      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       	          hff�?:ɨ��?            �@@�       �                   a@@4և���?
             ,@������������������������       �                     (@�       �                    @B@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?�\��N��?             3@�       �                    �K@�<ݚ�?             "@������������������������       �                     @�       �                    b@���Q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    �N@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @G@�z�G��?	             $@������������������������       �                     @�       �       	          ����?      �?             @������������������������       �                      @�       �       	          `ff@      �?             @������������������������       �                      @�       �                   �_@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                   �_@Xޒ�ZL�?           Py@�       �       	          ����?nM`����?8             W@�       �                    �?��v����?*            �P@�       �                   �b@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    @O@X��Oԣ�?'             O@�       �                    �E@ 	��p�?#             M@�       �                   �]@"pc�
�?             &@������������������������       �                      @�       �                   �Z@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?`�q�0ܴ?            �G@�       �                   �S@�(\����?             D@�       �                   �X@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                    �B@�       �       	             �?؇���X�?             @������������������������       �                     @������������������������       �                     �?�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     9@�       �       	          ����?���ס�?�            �s@�       �                    �?���5��?�            �q@�       �                   �j@�̚��?%            �N@�       �                   �f@���Q��?             $@�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?������?             �I@�       �                    �G@���@M^�?             ?@�       �                   �o@z�G�z�?             @������������������������       �                      @�       �                    �?�q�q�?             @�       �                    @F@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                   �c@�	j*D�?             :@�       �                   d@��<b���?             7@�       �                    �N@$�q-�?             *@������������������������       �                     $@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                     N@���Q��?             $@�       �                   `b@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     4@�       �                    I@����>��?�             l@�       �                     F@�q�q�?             (@������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @�       �       	          ���ٿz�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                   �c@ �h�7W�?�            �j@������������������������       �        D            @[@�       �                    �?\�t��Y�?H            �Y@�       �                    @I@��S���?             .@�       �                   �b@      �?              @������������������������       �                     @������������������������       �                      @�       �                    _@؇���X�?             @�       �                   0d@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �O@���7�?<             V@�       �                    @ ��N8�?:             U@������������������������       �        6             T@�       �                    �G@      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �d@      �?             @������������������������       �                     @������������������������       �                     �?�       �                   pb@d}h���?             <@�       �                    h@8�Z$���?             :@������������������������       �                     *@�       �                    �?�	j*D�?
             *@�       �                   `i@"pc�
�?	             &@������������������������       �                     �?�       �                    �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@������������������������       �                      @������������������������       �                      @�t�bh�h(h+K ��h-��R�(KK�KK��h_�B�        y@     0�@     �U@     �z@      U@     �z@     �I@     �x@             @X@     �I@     �r@       @      @      @       @               @      @              �?      @      �?                      @     �E@     @r@      6@      J@      ,@      @      (@       @              �?      (@      �?      @      �?      �?      �?      �?                      �?      @              @               @      @              @       @               @     �F@      @     �F@      @       @       @              �?       @      �?                       @      @     �E@      @      :@              &@      @      .@      @      @      �?               @      @               @       @      @              @       @                      "@              1@       @              5@      n@      @      0@       @      ,@              @       @       @      �?      �?      �?                      �?      �?      @      �?       @      �?      �?      �?                      �?              �?              @      @       @               @      @              .@      l@      "@      M@      �?      5@              2@      �?      @              @      �?               @     �B@       @      �?              �?       @              @      B@      �?      @@      �?       @              @      �?       @               @      �?                      8@      @      @              @      @              @     �d@       @     @Z@      �?     @W@      �?      5@              .@      �?      @      �?      �?              �?      �?                      @              R@      �?      (@              (@      �?              @     �N@      @      2@       @      @       @                      @       @      .@      �?      .@      �?                      .@      �?                     �E@     �@@      @@      7@      "@      7@      @      .@               @      @              @       @      @       @       @      �?      �?      �?                      �?      @      �?      @                      �?              �?              @      $@      7@      �?      *@              (@      �?      �?              �?      �?              "@      $@       @      @              @       @      @       @      �?      �?              �?      �?      �?                      �?               @      @      @      @              @      @               @      @      �?       @              �?      �?              �?      �?               @             �s@     �V@      M@      A@      M@      "@      @       @      @                       @     �K@      @      K@      @      "@       @       @              �?       @               @      �?             �F@       @     �C@      �?       @      �?              �?       @             �B@              @      �?      @                      �?      �?      @              @      �?                      9@      p@     �L@     @o@     �A@     �E@      2@      @      @      �?      @              @      �?              @             �C@      (@      3@      (@      �?      @               @      �?       @      �?      �?              �?      �?                      �?      2@       @      2@      @      (@      �?      $@               @      �?              �?       @              @      @      @      �?      @                      �?              @              @      4@             �i@      1@      @      @              @      @      �?      @              @      �?              �?      @              i@      (@     @[@             �V@      (@      @       @      @       @      @                       @      �?      @      �?      �?              �?      �?                      @      U@      @     �T@      �?      T@              @      �?       @              �?      �?      �?                      �?      �?      @              @      �?              @      6@      @      6@              *@      @      "@       @      "@      �?              �?      "@      �?                      "@       @               @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJe�MohG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvM3hwh(h+K ��h-��R�(KM3��h~�B(C         �                    @K@������?W           ��@       a                    �?    ��?B            �@       6                    �?������?�            @o@       )                    �?�n\�GZ�?K            �]@                          l@l��[B��?7            �U@                            E@�	j*D�?            �C@                           @D@�C��2(�?             &@������������������������       �                     @	       
                    ^@r�q��?             @������������������������       �                     �?������������������������       �                     @                           �?��>4և�?             <@              	             �?$��m��?             :@              
             �?X�<ݚ�?             2@������������������������       �                     @                           ]@���!pc�?             &@                           �E@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @                          �e@      �?              @                          `T@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @       (                    @J@      �?             H@                           �?�K��&�?            �E@������������������������       �                     @       '                    �H@P����?             C@       &       	          ����?<ݚ)�?             B@        %       
             �?r٣����?            �@@!       $                   (s@�q�q�?             (@"       #                   r@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     5@������������������������       �                     @������������������������       �                      @������������������������       �                     @*       +                    @I@      �?             @@������������������������       �        	             .@,       3                   ``@������?             1@-       .                    �?؇���X�?             ,@������������������������       �                     �?/       0                   �`@$�q-�?             *@������������������������       �                     @1       2       	          ����?r�q��?             @������������������������       �                     @������������������������       �                     �?4       5       
             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @7       8                   �U@���A���?I            ``@������������������������       �                     @9       Z       
             �? ��P0�?H            �_@:       Q                    �?@��xQ�??            �\@;       N                   �b@�8��8N�?6             X@<       E                    �?0�>���?3            �V@=       >                    �G@�θ�?             *@������������������������       �                     @?       @                   �k@�q�q�?             "@������������������������       �                     @A       B                   �p@���Q��?             @������������������������       �                      @C       D                   �s@�q�q�?             @������������������������       �                      @������������������������       �                     �?F       K                   pb@ ���J��?-            �S@G       H                   �_@`׀�:M�?+            �R@������������������������       �                     G@I       J                   pb@h�����?             <@������������������������       �                     ;@������������������������       �                     �?L       M                    �?      �?             @������������������������       �                     �?������������������������       �                     @O       P                    @E@���Q��?             @������������������������       �                     @������������������������       �                      @R       U                    @G@�<ݚ�?	             2@S       T                   �`@���Q��?             @������������������������       �                      @������������������������       �                     @V       Y                   �]@$�q-�?             *@W       X       	              @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @[       `                    @J@�n_Y�K�?	             *@\       _                   �`@z�G�z�?             $@]       ^                    @H@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @b       u       	          ����?��Eo5�?�            `p@c       n       
             �?��x��?�            @i@d       m       	          ����?�G�z��?             D@e       l                   0a@��<b���?             7@f       g                    @E@�q�q�?             .@������������������������       �                     @h       k                    �?�C��2(�?             &@i       j                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     1@o       t                   c@ A��� �?t            @d@p       s                    �? ����?1            @P@q       r                   �b@�h����?+             L@������������������������       �        *            �K@������������������������       �                     �?������������������������       �                     "@������������������������       �        C            @X@v       {                    �?*;L]n�?&             N@w       z       	          ����?�8��8��?	             (@x       y                   �b@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@|       �       
             �?�q���?             H@}       �                   �b@p�ݯ��?             C@~                          �i@�C��2(�?             6@������������������������       �                     *@�       �                   �l@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�       �       	             �?      �?             0@������������������������       �                     "@�       �                   (p@և���X�?             @�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    `@ףp=
�?             $@�       �                    �?z�G�z�?             @������������������������       �                      @�       �                   `d@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	          ����?x��ǃ�?           `y@�       �                   @E@��1���?n            �c@�       �                   �\@��-�=��?            �C@������������������������       �                     9@�       �       
             �?����X�?             ,@������������������������       �                     @�       �                    �?և���X�?             @�       �                    �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                    �?�0�w�?T            �]@�       �                   @b@H~��D
�?@            �W@�       �                   @e@z���=��?3            @S@�       �                   0r@�G�V�e�?-             Q@�       �                   �]@�j��b�?&            �M@�       �                     L@����X�?             @������������������������       �                      @������������������������       �                     @�       �                    �?$�q-�?"             J@�       �                    �L@"pc�
�?             &@�       �                    `@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       
             �?�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                    �Q@������?            �D@�       �                   Pa@�(\����?             D@������������������������       �                     5@�       �                    �?�}�+r��?             3@������������������������       �        
             0@�       �                   �h@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�       �                    `@�q�q�?             "@������������������������       �                     @�       �                    @      �?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    �?X�<ݚ�?             "@�       �                    �?z�G�z�?             @�       �                   f@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?X�<ݚ�?             2@�       �                    �N@����X�?
             ,@�       �                    �?���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    @�����H�?             "@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                    �N@      �?             8@�       �                    ]@      �?             0@�       �       
             �?r�q��?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �M@�z�G��?	             $@�       �                   Pd@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     @������������������������       �                     �?�       �                    �?�חF�P�?�             o@�       �                   �f@��S���?             >@������������������������       �                     @�       �                   Pd@� �	��?             9@�       �                    �?���|���?             6@�       �       
             �?������?             1@�       �                    �?X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @�       �                   �`@z�G�z�?             @�       �                   �q@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�                         �`@������?�            @k@�       �                    �?"pc�
�?8             V@�       �                   Xy@�8��8��?&             N@�       �       
             �? ,��-�?%            �M@�       �                    \@�&=�w��?!            �J@�       �                    @M@8�Z$���?             *@�       �                   �Y@���Q��?             @������������������������       �                     �?�       �                   �`@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     D@�       �                   �]@�q�q�?             @������������������������       �                      @�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     �?                          c@��>4և�?             <@      
      	          `ff�?��.k���?             1@                         �?�	j*D�?             *@������������������������       �                     �?      	                  �_@      �?             (@                        Pr@      �?              @                         �O@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @                         �?"pc�
�?             &@                         �L@ףp=
�?             $@                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?      0                   �R@$�q-�?W            @`@      '      
             �?     ��?U             `@                         �?�8���?K             ]@                         �?؇���X�?             <@                         @����X�?
             ,@                        �]@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@                        �a@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     ,@                          �?`���i��?9             V@������������������������       �        /             R@!      &                  �n@      �?
             0@"      %                  pm@z�G�z�?             $@#      $                  �e@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @(      /                  �p@      �?
             (@)      .                   e@"pc�
�?	             &@*      +      	          ��� @ףp=
�?             $@������������������������       �                      @,      -                   o@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?1      2                  �b@      �?              @������������������������       �                     �?������������������������       �                     �?�t�bh�h(h+K ��h-��R�(KM3KK��h_�B0       �y@     �@     �q@     �l@     �P@      g@      G@     @R@      E@     �F@      (@      ;@      �?      $@              @      �?      @      �?                      @      &@      1@      "@      1@       @      $@              @       @      @       @      @       @                      @      @              �?      @      �?       @               @      �?                      @       @              >@      2@      9@      2@              @      9@      *@      9@      &@      9@       @      @       @      @      @              @      @                      @      5@                      @               @      @              @      <@              .@      @      *@       @      (@      �?              �?      (@              @      �?      @              @      �?               @      �?              �?       @              4@     �[@      @              0@     �[@      &@     �Y@      @     @V@      @     �U@      @      $@              @      @      @              @      @       @       @              �?       @               @      �?               @      S@      �?     @R@              G@      �?      ;@              ;@      �?              �?      @      �?                      @       @      @              @       @              @      ,@      @       @               @      @              �?      (@      �?      @              @      �?                       @      @       @       @       @       @      @       @                      @              @      @              k@     �F@     �f@      3@      6@      2@      @      2@      @      $@      @              �?      $@      �?       @      �?                       @               @               @      1@              d@      �?      P@      �?     �K@      �?     �K@                      �?      "@             @X@              A@      :@      &@      �?      �?      �?      �?                      �?      $@              7@      9@      ,@      8@       @      4@              *@       @      @       @                      @      (@      @      "@              @      @      @      �?      @                      �?              @      "@      �?      @      �?       @               @      �?       @                      �?      @             �_@     pq@     �U@     �Q@      @     �A@              9@      @      $@              @      @      @      @       @      @                       @              �?     �T@      B@     �R@      5@      P@      *@     �M@      "@     �J@      @      @       @               @      @              H@      @      "@       @      �?      �?              �?      �?               @      �?              �?       @             �C@       @     �C@      �?      5@              2@      �?      0@               @      �?       @                      �?              �?      @      @      @              @      @      @      �?              �?      @                       @      @      @      �?      @      �?       @               @      �?                       @      @              $@       @      $@      @       @      @              @       @               @      �?      �?      �?      �?                      �?      @                      @      "@      .@       @       @      @      �?      �?      �?      �?                      �?      @              @      @      @      @              @      @                      @      �?      @              @      �?              D@      j@      ,@      0@              @      ,@      &@      ,@       @      *@      @      @      @              @      @               @              �?      @      �?      �?              �?      �?                      @              @      :@      h@      0@      R@      @     �K@      @     �K@       @     �I@       @      &@       @      @              �?       @       @       @                       @               @              D@       @      @               @       @       @       @                       @      �?              &@      1@      "@       @      "@      @              �?      "@      @      @      @      @      �?              �?      @                       @      @                      @       @      "@      �?      "@      �?       @      �?                       @              @      �?              $@      ^@      "@     �]@      @     �[@      @      8@      @      $@      �?      "@      �?                      "@      @      �?              �?      @                      ,@       @     �U@              R@       @      ,@       @       @      �?       @               @      �?              �?                      @      @      "@       @      "@      �?      "@               @      �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��lhG        hNhG        hEKhFKhGh(h+K ��h-��R�(KK��h_�C              �?�t�bhShdhNC       ���R�hhKhihlKh(h+K ��h-��R�(KK��hN�C       �t�bK��R�}�(hKhvK�hwh(h+K ��h-��R�(KK���h~�B�7         �       
             �?�HK��x�?>           ��@       W                    �?8z^����?F           Ѐ@                          �`@�P+SS�?~            `j@              
             �?l�b�G��?#            �L@������������������������       �                     @                           �?HP�s��?             I@                          c@      �?              @������������������������       �                     @	       
                    �?      �?             @������������������������       �                     �?������������������������       �                     @                          �^@�Ń��̧?             E@                           �?�IєX�?             1@������������������������       �        	             .@                          �Z@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     9@       0                    �?$;hB��?[            @c@       +                    �?��h!��?$            �L@                          @]@(���@��?            �G@������������������������       �                     &@                           �?�q�q�?             B@                           �M@�q�q�?             "@������������������������       �                     @                            O@���Q��?             @������������������������       �                     @������������������������       �                      @       $                    �K@�q�q�?             ;@       #                   �d@@�0�!��?	             1@                           �q@      �?             0@������������������������       �                     $@!       "                    @G@�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?%       *                   �d@���Q��?             $@&       )                    b@      �?              @'       (       	             �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @,       -       	          433�?ףp=
�?             $@������������������������       �                     @.       /                   �S@      �?             @������������������������       �                     �?������������������������       �                     @1       V                   f@����l�?7            @X@2       I                   Hp@��S���?3            �V@3       4                   g@��h!��?             �L@������������������������       �                     @5       :                    �?`�Q��?             I@6       9       	          @33�?�LQ�1	�?             7@7       8                    �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     .@;       @                    �L@|��?���?             ;@<       =       	          ����?z�G�z�?             $@������������������������       �                     �?>       ?                   �g@�����H�?             "@������������������������       �                     �?������������������������       �                      @A       B       	          pff�?ҳ�wY;�?             1@������������������������       �                     @C       D                    `@8�Z$���?             *@������������������������       �                     @E       F       	          `ff�?�<ݚ�?             "@������������������������       �                     @G       H                    �N@���Q��?             @������������������������       �                     @������������������������       �                      @J       U                   �@�'�`d�?            �@@K       R                    �?�r����?             >@L       M                   �p@      �?             @������������������������       �                     �?N       Q       	          `ff�?���Q��?             @O       P                    �N@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @S       T       	          ���@ �q�q�?             8@������������������������       �                     7@������������������������       �                     �?������������������������       �                     @������������������������       �                     @X       �                   �b@��<nd�?�            pt@Y       �                    @�IєX�?�             s@Z       }                   P`@����?�             s@[       l                    �?���	���?O             a@\       ]       
             �?P���Q�?9             Y@������������������������       �        
             1@^       a                    �? ,U,?��?/            �T@_       `                   @_@�q�q�?             @������������������������       �                      @������������������������       �                     �?b       i                    `P@x�G�z�?-             T@c       d                    `@�k~X��?)             R@������������������������       �                     K@e       f                   �s@�X�<ݺ?             2@������������������������       �        
             0@g       h                   �|@      �?              @������������������������       �                     �?������������������������       �                     �?j       k                    Y@      �?              @������������������������       �                      @������������������������       �                     @m       |       	             @���@��?            �B@n       q                    �G@b�h�d.�?            �A@o       p                    �F@���Q��?             @������������������������       �                     @������������������������       �                      @r       {       	          ����?�r����?             >@s       t       	             �?�q�q�?	             (@������������������������       �                     @u       z                    �M@      �?              @v       y                   �X@�q�q�?             @w       x                    @K@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �        
             2@������������������������       �                      @~                          �j@ d��?k            �d@������������������������       �        ,            @Q@�       �                    �R@@9G��??            �X@�       �       	          ����?      �?=             X@�       �                    �?�����H�?             2@�       �                   �`@r�q��?             (@�       �                   �_@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                   k@�(�Tw�?0            �S@�       �                   �a@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        .             S@�       �       
             �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �[@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   �q@և���X�?             5@�       �       	          033�?     ��?
             0@�       �                   �b@      �?              @������������������������       �                     @������������������������       �                     �?�       �                   �p@      �?              @�       �                    c@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   @E@>���$��?�            �w@�       �                   `@�+e�X�?              I@�       �                   a@���}<S�?             7@������������������������       �        
             1@�       �                   �]@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                   �b@��}*_��?             ;@�       �                    �?��+7��?             7@�       �                     L@�q�q�?             "@�       �                   �\@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     ,@������������������������       �                     @�       �       	          033@�r����?�            �t@�       �                    �?����ր�?�            @t@�       �                    �?      �?&             L@�       �                    �?R���Q�?             4@�       �                   ps@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     *@�       �                   d@      �?             B@�       �                     I@�X����?             6@������������������������       �                     (@�       �                    @O@�z�G��?             $@������������������������       �                     @�       �       	          `ff @      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?d}h���?             ,@�       �                   Pq@�θ�?
             *@�       �                    �?ףp=
�?             $@�       �                    �?؇���X�?             @������������������������       �                      @�       �                    @L@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                   Pe@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �       	             �?��	��j�?�            �p@�       �                    �I@ $i���?�            �m@�       �                   @[@�|�l�?S             a@�       �                   �b@��S�ۿ?
             .@������������������������       �                     @�       �                   �c@      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �        I            @^@�       �                    @J@�:�]��?E            �Y@�       �                   pl@������?             .@������������������������       �                     @�       �                   p@      �?              @������������������������       �                     @������������������������       �                     @�       �                    �?`��F:u�?:            �U@�       �                    �?r�q��?             2@������������������������       �                     @�       �                    �?      �?
             (@�       �                   �h@�z�G��?	             $@������������������������       �                     @�       �                    �M@���Q��?             @�       �       	          ����?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                   �a@@	tbA@�?-            @Q@������������������������       �                    �B@�       �                   �a@      �?             @@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     =@�       �                    �?������?             >@�       �                    k@r�q��?             8@�       �                     I@�q�q�?             "@������������������������       �                     @�       �       	          ����?      �?             @������������������������       �                     @������������������������       �                     @�       �       	          ����?��S�ۿ?             .@������������������������       �                     $@�       �                   �`@z�G�z�?             @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     M@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�t�b�'      h�h(h+K ��h-��R�(KK�KK��h_�B�        y@     0�@     �Y@     @{@     �R@      a@      @     �J@              @      @      G@      @      @              @      @      �?              �?      @              �?     �D@      �?      0@              .@      �?      �?      �?                      �?              9@     �Q@     �T@      0@     �D@      .@      @@              &@      .@      5@      @      @      @               @      @              @       @              "@      2@      @      ,@       @      ,@              $@       @      @              @       @              �?              @      @      @       @      �?       @      �?                       @      @                       @      �?      "@              @      �?      @      �?                      @     �K@      E@      H@      E@     �D@      0@      @              A@      0@      4@      @      @      @              @      @              .@              ,@      *@       @       @              �?       @      �?              �?       @              @      &@      @               @      &@              @       @      @              @       @      @              @       @              @      :@      @      :@      @      @              �?      @       @      �?       @               @      �?               @              �?      7@              7@      �?              @              @              ;@     �r@      2@      r@      1@     �q@      *@      _@      @     �W@              1@      @     �S@       @      �?       @                      �?      @     @S@      �?     �Q@              K@      �?      1@              0@      �?      �?      �?                      �?       @      @       @                      @       @      =@      @      =@       @      @              @       @              @      :@      @       @              @      @      @       @      @       @      �?              �?       @                      @       @                      2@       @              @     `d@             @Q@      @     �W@      @     @W@       @      0@       @      $@       @       @               @       @                       @              @      �?     @S@      �?      �?      �?                      �?              S@      �?      �?      �?                      �?      �?      �?      �?                      �?      "@      (@      "@      @      @      �?      @                      �?       @      @      �?      @      �?                      @      �?                      @     �r@     �T@      (@      C@       @      5@              1@       @      @       @                      @      $@      1@      @      1@      @      @       @      @       @                      @      @                      ,@      @             �q@      F@     �q@      C@     �A@      5@      1@      @      @      @      @                      @      *@              2@      2@      @      .@              (@      @      @      @              �?      @              @      �?              &@      @      $@      @      "@      �?      @      �?       @              @      �?      @                      �?      @              �?       @      �?                       @      �?             `o@      1@     �l@      "@     �`@      �?      ,@      �?      @              @      �?              �?      @             @^@             �W@       @      &@      @      @              @      @              @      @             �T@      @      .@      @      @              "@      @      @      @      @               @      @       @      �?       @                      �?               @       @              Q@      �?     �B@              ?@      �?       @      �?              �?       @              =@              6@       @      4@      @      @      @      @              @      @              @      @              ,@      �?      $@              @      �?      @              �?      �?      �?                      �?       @      @       @                      @              @�t�bubhhubehhub.